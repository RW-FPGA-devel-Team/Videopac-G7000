-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d5",
     9 => x"b4080b0b",
    10 => x"80d5b808",
    11 => x"0b0b80d5",
    12 => x"bc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d5bc0c0b",
    16 => x"0b80d5b8",
    17 => x"0c0b0b80",
    18 => x"d5b40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b80cad4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d5b470",
    57 => x"80dfec27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c5197c5",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d5",
    65 => x"c40c9f0b",
    66 => x"80d5c80c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d5c808ff",
    70 => x"0580d5c8",
    71 => x"0c80d5c8",
    72 => x"088025e8",
    73 => x"3880d5c4",
    74 => x"08ff0580",
    75 => x"d5c40c80",
    76 => x"d5c40880",
    77 => x"25d03880",
    78 => x"0b80d5c8",
    79 => x"0c800b80",
    80 => x"d5c40c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d5c408",
   100 => x"25913882",
   101 => x"c82d80d5",
   102 => x"c408ff05",
   103 => x"80d5c40c",
   104 => x"838a0480",
   105 => x"d5c40880",
   106 => x"d5c80853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d5c408",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d5c80881",
   116 => x"0580d5c8",
   117 => x"0c80d5c8",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d5c8",
   121 => x"0c80d5c4",
   122 => x"08810580",
   123 => x"d5c40c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d5",
   128 => x"c8088105",
   129 => x"80d5c80c",
   130 => x"80d5c808",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d5c8",
   134 => x"0c80d5c4",
   135 => x"08810580",
   136 => x"d5c40c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d5cc0cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d5cc0c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d5",
   177 => x"cc088407",
   178 => x"80d5cc0c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5485bc74",
   182 => x"258f3882",
   183 => x"0b0b0b80",
   184 => x"d0800c80",
   185 => x"d05385f3",
   186 => x"04810b0b",
   187 => x"0b80d080",
   188 => x"0cbc530b",
   189 => x"0b80d080",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0cfc0875",
   193 => x"7531ffb0",
   194 => x"05ff1371",
   195 => x"712cff94",
   196 => x"1a709f2a",
   197 => x"1170812c",
   198 => x"80d5cc08",
   199 => x"52545153",
   200 => x"57535152",
   201 => x"5276802e",
   202 => x"85387081",
   203 => x"075170f6",
   204 => x"940c7209",
   205 => x"8105f680",
   206 => x"0c710981",
   207 => x"05f6840c",
   208 => x"0294050d",
   209 => x"0402f405",
   210 => x"0d745372",
   211 => x"70810554",
   212 => x"80f52d52",
   213 => x"71802e89",
   214 => x"38715183",
   215 => x"842d86cb",
   216 => x"04810b80",
   217 => x"d5b40c02",
   218 => x"8c050d04",
   219 => x"02fc050d",
   220 => x"81808051",
   221 => x"c0115170",
   222 => x"fb380284",
   223 => x"050d0402",
   224 => x"fc050dec",
   225 => x"5183710c",
   226 => x"86ec2d82",
   227 => x"710c0284",
   228 => x"050d0486",
   229 => x"ec2d86ec",
   230 => x"2d86ec2d",
   231 => x"86ec2d86",
   232 => x"ec2d86ec",
   233 => x"2d86ec2d",
   234 => x"86ec2d86",
   235 => x"ec2d86ec",
   236 => x"2d86ec2d",
   237 => x"86ec2d86",
   238 => x"ec2d86ec",
   239 => x"2d86ec2d",
   240 => x"86ec2d86",
   241 => x"ec2d86ec",
   242 => x"2d86ec2d",
   243 => x"86ec2d86",
   244 => x"ec2d86ec",
   245 => x"2d86ec2d",
   246 => x"86ec2d86",
   247 => x"ec2d86ec",
   248 => x"2d86ec2d",
   249 => x"86ec2d86",
   250 => x"ec2d86ec",
   251 => x"2d86ec2d",
   252 => x"86ec2d86",
   253 => x"ec2d86ec",
   254 => x"2d86ec2d",
   255 => x"86ec2d86",
   256 => x"ec2d86ec",
   257 => x"2d86ec2d",
   258 => x"86ec2d86",
   259 => x"ec2d86ec",
   260 => x"2d86ec2d",
   261 => x"86ec2d86",
   262 => x"ec2d86ec",
   263 => x"2d86ec2d",
   264 => x"86ec2d86",
   265 => x"ec2d86ec",
   266 => x"2d86ec2d",
   267 => x"86ec2d86",
   268 => x"ec2d86ec",
   269 => x"2d86ec2d",
   270 => x"86ec2d86",
   271 => x"ec2d86ec",
   272 => x"2d86ec2d",
   273 => x"86ec2d86",
   274 => x"ec2d86ec",
   275 => x"2d86ec2d",
   276 => x"86ec2d86",
   277 => x"ec2d86ec",
   278 => x"2d86ec2d",
   279 => x"86ec2d86",
   280 => x"ec2d86ec",
   281 => x"2d86ec2d",
   282 => x"86ec2d86",
   283 => x"ec2d86ec",
   284 => x"2d86ec2d",
   285 => x"86ec2d86",
   286 => x"ec2d86ec",
   287 => x"2d86ec2d",
   288 => x"86ec2d86",
   289 => x"ec2d86ec",
   290 => x"2d86ec2d",
   291 => x"86ec2d86",
   292 => x"ec2d86ec",
   293 => x"2d86ec2d",
   294 => x"86ec2d86",
   295 => x"ec2d86ec",
   296 => x"2d86ec2d",
   297 => x"86ec2d86",
   298 => x"ec2d86ec",
   299 => x"2d86ec2d",
   300 => x"86ec2d86",
   301 => x"ec2d86ec",
   302 => x"2d86ec2d",
   303 => x"86ec2d86",
   304 => x"ec2d86ec",
   305 => x"2d86ec2d",
   306 => x"86ec2d86",
   307 => x"ec2d86ec",
   308 => x"2d86ec2d",
   309 => x"86ec2d86",
   310 => x"ec2d86ec",
   311 => x"2d86ec2d",
   312 => x"86ec2d86",
   313 => x"ec2d86ec",
   314 => x"2d86ec2d",
   315 => x"86ec2d86",
   316 => x"ec2d86ec",
   317 => x"2d86ec2d",
   318 => x"86ec2d86",
   319 => x"ec2d86ec",
   320 => x"2d86ec2d",
   321 => x"86ec2d86",
   322 => x"ec2d86ec",
   323 => x"2d86ec2d",
   324 => x"86ec2d86",
   325 => x"ec2d86ec",
   326 => x"2d86ec2d",
   327 => x"86ec2d86",
   328 => x"ec2d86ec",
   329 => x"2d86ec2d",
   330 => x"86ec2d86",
   331 => x"ec2d86ec",
   332 => x"2d86ec2d",
   333 => x"86ec2d86",
   334 => x"ec2d86ec",
   335 => x"2d86ec2d",
   336 => x"86ec2d86",
   337 => x"ec2d86ec",
   338 => x"2d86ec2d",
   339 => x"86ec2d86",
   340 => x"ec2d86ec",
   341 => x"2d86ec2d",
   342 => x"86ec2d86",
   343 => x"ec2d86ec",
   344 => x"2d86ec2d",
   345 => x"86ec2d86",
   346 => x"ec2d86ec",
   347 => x"2d86ec2d",
   348 => x"86ec2d86",
   349 => x"ec2d86ec",
   350 => x"2d86ec2d",
   351 => x"86ec2d86",
   352 => x"ec2d86ec",
   353 => x"2d86ec2d",
   354 => x"86ec2d86",
   355 => x"ec2d86ec",
   356 => x"2d86ec2d",
   357 => x"86ec2d86",
   358 => x"ec2d86ec",
   359 => x"2d86ec2d",
   360 => x"86ec2d86",
   361 => x"ec2d86ec",
   362 => x"2d86ec2d",
   363 => x"86ec2d86",
   364 => x"ec2d86ec",
   365 => x"2d86ec2d",
   366 => x"86ec2d86",
   367 => x"ec2d86ec",
   368 => x"2d86ec2d",
   369 => x"86ec2d86",
   370 => x"ec2d86ec",
   371 => x"2d86ec2d",
   372 => x"86ec2d86",
   373 => x"ec2d86ec",
   374 => x"2d86ec2d",
   375 => x"86ec2d86",
   376 => x"ec2d86ec",
   377 => x"2d86ec2d",
   378 => x"86ec2d86",
   379 => x"ec2d86ec",
   380 => x"2d86ec2d",
   381 => x"86ec2d86",
   382 => x"ec2d86ec",
   383 => x"2d86ec2d",
   384 => x"86ec2d86",
   385 => x"ec2d86ec",
   386 => x"2d86ec2d",
   387 => x"86ec2d86",
   388 => x"ec2d86ec",
   389 => x"2d86ec2d",
   390 => x"86ec2d86",
   391 => x"ec2d86ec",
   392 => x"2d86ec2d",
   393 => x"86ec2d86",
   394 => x"ec2d86ec",
   395 => x"2d86ec2d",
   396 => x"86ec2d86",
   397 => x"ec2d86ec",
   398 => x"2d86ec2d",
   399 => x"86ec2d86",
   400 => x"ec2d86ec",
   401 => x"2d86ec2d",
   402 => x"86ec2d86",
   403 => x"ec2d86ec",
   404 => x"2d86ec2d",
   405 => x"86ec2d86",
   406 => x"ec2d86ec",
   407 => x"2d86ec2d",
   408 => x"86ec2d86",
   409 => x"ec2d86ec",
   410 => x"2d86ec2d",
   411 => x"86ec2d86",
   412 => x"ec2d86ec",
   413 => x"2d86ec2d",
   414 => x"86ec2d86",
   415 => x"ec2d86ec",
   416 => x"2d86ec2d",
   417 => x"86ec2d86",
   418 => x"ec2d86ec",
   419 => x"2d86ec2d",
   420 => x"86ec2d86",
   421 => x"ec2d86ec",
   422 => x"2d86ec2d",
   423 => x"86ec2d86",
   424 => x"ec2d86ec",
   425 => x"2d86ec2d",
   426 => x"86ec2d86",
   427 => x"ec2d86ec",
   428 => x"2d86ec2d",
   429 => x"86ec2d86",
   430 => x"ec2d86ec",
   431 => x"2d86ec2d",
   432 => x"86ec2d86",
   433 => x"ec2d86ec",
   434 => x"2d86ec2d",
   435 => x"86ec2d86",
   436 => x"ec2d86ec",
   437 => x"2d86ec2d",
   438 => x"86ec2d86",
   439 => x"ec2d86ec",
   440 => x"2d86ec2d",
   441 => x"86ec2d86",
   442 => x"ec2d86ec",
   443 => x"2d86ec2d",
   444 => x"86ec2d86",
   445 => x"ec2d86ec",
   446 => x"2d86ec2d",
   447 => x"86ec2d86",
   448 => x"ec2d86ec",
   449 => x"2d86ec2d",
   450 => x"86ec2d86",
   451 => x"ec2d86ec",
   452 => x"2d86ec2d",
   453 => x"86ec2d86",
   454 => x"ec2d86ec",
   455 => x"2d86ec2d",
   456 => x"86ec2d86",
   457 => x"ec2d86ec",
   458 => x"2d86ec2d",
   459 => x"86ec2d86",
   460 => x"ec2d86ec",
   461 => x"2d86ec2d",
   462 => x"86ec2d86",
   463 => x"ec2d86ec",
   464 => x"2d86ec2d",
   465 => x"86ec2d86",
   466 => x"ec2d86ec",
   467 => x"2d86ec2d",
   468 => x"86ec2d86",
   469 => x"ec2d86ec",
   470 => x"2d86ec2d",
   471 => x"86ec2d86",
   472 => x"ec2d86ec",
   473 => x"2d86ec2d",
   474 => x"86ec2d86",
   475 => x"ec2d86ec",
   476 => x"2d86ec2d",
   477 => x"86ec2d86",
   478 => x"ec2d86ec",
   479 => x"2d86ec2d",
   480 => x"86ec2d86",
   481 => x"ec2d86ec",
   482 => x"2d86ec2d",
   483 => x"86ec2d86",
   484 => x"ec2d86ec",
   485 => x"2d86ec2d",
   486 => x"86ec2d86",
   487 => x"ec2d86ec",
   488 => x"2d86ec2d",
   489 => x"86ec2d86",
   490 => x"ec2d86ec",
   491 => x"2d86ec2d",
   492 => x"86ec2d86",
   493 => x"ec2d86ec",
   494 => x"2d86ec2d",
   495 => x"86ec2d86",
   496 => x"ec2d86ec",
   497 => x"2d86ec2d",
   498 => x"86ec2d86",
   499 => x"ec2d86ec",
   500 => x"2d86ec2d",
   501 => x"86ec2d86",
   502 => x"ec2d86ec",
   503 => x"2d86ec2d",
   504 => x"86ec2d86",
   505 => x"ec2d86ec",
   506 => x"2d86ec2d",
   507 => x"86ec2d86",
   508 => x"ec2d86ec",
   509 => x"2d86ec2d",
   510 => x"86ec2d86",
   511 => x"ec2d86ec",
   512 => x"2d86ec2d",
   513 => x"86ec2d86",
   514 => x"ec2d86ec",
   515 => x"2d86ec2d",
   516 => x"86ec2d86",
   517 => x"ec2d86ec",
   518 => x"2d86ec2d",
   519 => x"86ec2d86",
   520 => x"ec2d86ec",
   521 => x"2d86ec2d",
   522 => x"86ec2d86",
   523 => x"ec2d86ec",
   524 => x"2d86ec2d",
   525 => x"86ec2d86",
   526 => x"ec2d86ec",
   527 => x"2d86ec2d",
   528 => x"86ec2d86",
   529 => x"ec2d86ec",
   530 => x"2d86ec2d",
   531 => x"86ec2d86",
   532 => x"ec2d86ec",
   533 => x"2d86ec2d",
   534 => x"86ec2d86",
   535 => x"ec2d86ec",
   536 => x"2d86ec2d",
   537 => x"86ec2d86",
   538 => x"ec2d86ec",
   539 => x"2d86ec2d",
   540 => x"86ec2d86",
   541 => x"ec2d86ec",
   542 => x"2d86ec2d",
   543 => x"86ec2d86",
   544 => x"ec2d86ec",
   545 => x"2d86ec2d",
   546 => x"86ec2d86",
   547 => x"ec2d86ec",
   548 => x"2d86ec2d",
   549 => x"86ec2d86",
   550 => x"ec2d86ec",
   551 => x"2d86ec2d",
   552 => x"86ec2d86",
   553 => x"ec2d86ec",
   554 => x"2d86ec2d",
   555 => x"86ec2d86",
   556 => x"ec2d86ec",
   557 => x"2d86ec2d",
   558 => x"86ec2d86",
   559 => x"ec2d86ec",
   560 => x"2d86ec2d",
   561 => x"86ec2d86",
   562 => x"ec2d86ec",
   563 => x"2d86ec2d",
   564 => x"86ec2d86",
   565 => x"ec2d86ec",
   566 => x"2d86ec2d",
   567 => x"86ec2d86",
   568 => x"ec2d86ec",
   569 => x"2d86ec2d",
   570 => x"86ec2d86",
   571 => x"ec2d86ec",
   572 => x"2d86ec2d",
   573 => x"86ec2d86",
   574 => x"ec2d86ec",
   575 => x"2d86ec2d",
   576 => x"86ec2d86",
   577 => x"ec2d86ec",
   578 => x"2d86ec2d",
   579 => x"86ec2d86",
   580 => x"ec2d86ec",
   581 => x"2d86ec2d",
   582 => x"86ec2d86",
   583 => x"ec2d86ec",
   584 => x"2d86ec2d",
   585 => x"86ec2d86",
   586 => x"ec2d86ec",
   587 => x"2d86ec2d",
   588 => x"86ec2d86",
   589 => x"ec2d86ec",
   590 => x"2d86ec2d",
   591 => x"86ec2d86",
   592 => x"ec2d86ec",
   593 => x"2d86ec2d",
   594 => x"86ec2d86",
   595 => x"ec2d86ec",
   596 => x"2d86ec2d",
   597 => x"86ec2d86",
   598 => x"ec2d86ec",
   599 => x"2d86ec2d",
   600 => x"86ec2d86",
   601 => x"ec2d86ec",
   602 => x"2d86ec2d",
   603 => x"86ec2d86",
   604 => x"ec2d86ec",
   605 => x"2d86ec2d",
   606 => x"86ec2d86",
   607 => x"ec2d86ec",
   608 => x"2d86ec2d",
   609 => x"86ec2d86",
   610 => x"ec2d86ec",
   611 => x"2d86ec2d",
   612 => x"86ec2d86",
   613 => x"ec2d86ec",
   614 => x"2d86ec2d",
   615 => x"86ec2d86",
   616 => x"ec2d86ec",
   617 => x"2d86ec2d",
   618 => x"86ec2d86",
   619 => x"ec2d86ec",
   620 => x"2d86ec2d",
   621 => x"86ec2d86",
   622 => x"ec2d86ec",
   623 => x"2d86ec2d",
   624 => x"86ec2d86",
   625 => x"ec2d86ec",
   626 => x"2d86ec2d",
   627 => x"86ec2d86",
   628 => x"ec2d86ec",
   629 => x"2d86ec2d",
   630 => x"86ec2d86",
   631 => x"ec2d86ec",
   632 => x"2d86ec2d",
   633 => x"86ec2d86",
   634 => x"ec2d86ec",
   635 => x"2d86ec2d",
   636 => x"86ec2d86",
   637 => x"ec2d86ec",
   638 => x"2d86ec2d",
   639 => x"86ec2d86",
   640 => x"ec2d86ec",
   641 => x"2d86ec2d",
   642 => x"86ec2d86",
   643 => x"ec2d86ec",
   644 => x"2d86ec2d",
   645 => x"86ec2d86",
   646 => x"ec2d86ec",
   647 => x"2d86ec2d",
   648 => x"86ec2d86",
   649 => x"ec2d86ec",
   650 => x"2d86ec2d",
   651 => x"86ec2d86",
   652 => x"ec2d86ec",
   653 => x"2d86ec2d",
   654 => x"86ec2d86",
   655 => x"ec2d86ec",
   656 => x"2d86ec2d",
   657 => x"86ec2d86",
   658 => x"ec2d86ec",
   659 => x"2d86ec2d",
   660 => x"86ec2d04",
   661 => x"0402dc05",
   662 => x"0d7a5580",
   663 => x"59840bec",
   664 => x"0c80d088",
   665 => x"085380d0",
   666 => x"8408812e",
   667 => x"0981068c",
   668 => x"38728280",
   669 => x"0780d088",
   670 => x"0c958704",
   671 => x"72828007",
   672 => x"82803280",
   673 => x"d0880c80",
   674 => x"d08808fc",
   675 => x"0c86ec2d",
   676 => x"745280d5",
   677 => x"d05180c0",
   678 => x"f62d80d5",
   679 => x"b408802e",
   680 => x"81c63880",
   681 => x"d5d40854",
   682 => x"80567385",
   683 => x"2e098106",
   684 => x"bb387451",
   685 => x"86c52d87",
   686 => x"932d8793",
   687 => x"2d87932d",
   688 => x"87932d87",
   689 => x"932d8793",
   690 => x"2d80d684",
   691 => x"08882a70",
   692 => x"81065153",
   693 => x"72762e88",
   694 => x"3880d1b4",
   695 => x"5195e404",
   696 => x"80d08c51",
   697 => x"a2982d81",
   698 => x"5397bb04",
   699 => x"73f80ca5",
   700 => x"0bec0c87",
   701 => x"932d840b",
   702 => x"ec0c75ff",
   703 => x"15575875",
   704 => x"802e8b38",
   705 => x"81187681",
   706 => x"2a575895",
   707 => x"ff04f718",
   708 => x"58815980",
   709 => x"742580d0",
   710 => x"38775275",
   711 => x"5184a82d",
   712 => x"80d6a452",
   713 => x"80d5d051",
   714 => x"80c3c82d",
   715 => x"80d5b408",
   716 => x"802e9b38",
   717 => x"80d6a457",
   718 => x"83fc5576",
   719 => x"70840558",
   720 => x"08e80cfc",
   721 => x"15557480",
   722 => x"25f13896",
   723 => x"d60480d5",
   724 => x"b4085984",
   725 => x"805480d5",
   726 => x"d05180c3",
   727 => x"982dfc80",
   728 => x"14811757",
   729 => x"54969304",
   730 => x"80d08408",
   731 => x"53728938",
   732 => x"725186ff",
   733 => x"2d978f04",
   734 => x"800b80d0",
   735 => x"840c80d0",
   736 => x"88088280",
   737 => x"07828032",
   738 => x"7080d088",
   739 => x"0cfc0c78",
   740 => x"802e9f38",
   741 => x"80d68408",
   742 => x"882a7081",
   743 => x"06515372",
   744 => x"802e8838",
   745 => x"80d1b451",
   746 => x"97b60480",
   747 => x"d08c5197",
   748 => x"b60480d2",
   749 => x"dc51a298",
   750 => x"2d785372",
   751 => x"80d5b40c",
   752 => x"02a4050d",
   753 => x"0402e805",
   754 => x"0d805186",
   755 => x"ff2d840b",
   756 => x"ec0c9fb0",
   757 => x"2d9bdb2d",
   758 => x"81f92d83",
   759 => x"539f932d",
   760 => x"8151858d",
   761 => x"2dff1353",
   762 => x"728025f1",
   763 => x"38840bec",
   764 => x"0c80ceb4",
   765 => x"5186c52d",
   766 => x"b7aa2d80",
   767 => x"d5b40880",
   768 => x"2e83c138",
   769 => x"810bec0c",
   770 => x"840bec0c",
   771 => x"80cae452",
   772 => x"80d5d051",
   773 => x"80c0f62d",
   774 => x"80d5b408",
   775 => x"802e80cc",
   776 => x"3880d6a4",
   777 => x"5280d5d0",
   778 => x"5180c3c8",
   779 => x"2d80d5b4",
   780 => x"08802eb8",
   781 => x"3880d6a4",
   782 => x"0b80f52d",
   783 => x"80d3e00c",
   784 => x"80d6a50b",
   785 => x"80f52d80",
   786 => x"d3e40c80",
   787 => x"d6a60b80",
   788 => x"f52d80d3",
   789 => x"e80c80d6",
   790 => x"a70b80f5",
   791 => x"2d80d3ec",
   792 => x"0c80d6a8",
   793 => x"0b80f52d",
   794 => x"80d3f00c",
   795 => x"80caf452",
   796 => x"80d5d051",
   797 => x"80c0f62d",
   798 => x"80d5b408",
   799 => x"802e80cc",
   800 => x"3880d6a4",
   801 => x"5280d5d0",
   802 => x"5180c3c8",
   803 => x"2d80d5b4",
   804 => x"08802eb8",
   805 => x"3880d6a4",
   806 => x"0b80f52d",
   807 => x"80d3cc0c",
   808 => x"80d6a50b",
   809 => x"80f52d80",
   810 => x"d3d00c80",
   811 => x"d6a60b80",
   812 => x"f52d80d3",
   813 => x"d40c80d6",
   814 => x"a70b80f5",
   815 => x"2d80d3d8",
   816 => x"0c80d6a8",
   817 => x"0b80f52d",
   818 => x"80d3dc0c",
   819 => x"94d55180",
   820 => x"cacc2d80",
   821 => x"d0880880",
   822 => x"d3c80c80",
   823 => x"d08808fc",
   824 => x"0c80d684",
   825 => x"08882a70",
   826 => x"81065153",
   827 => x"72802e88",
   828 => x"3880d1b4",
   829 => x"5199fc04",
   830 => x"80d08c51",
   831 => x"a2982d86",
   832 => x"0b80d698",
   833 => x"0c9fe92d",
   834 => x"9be72da2",
   835 => x"ab2d80d5",
   836 => x"b40880d6",
   837 => x"8408882a",
   838 => x"70810651",
   839 => x"54557280",
   840 => x"2ead3880",
   841 => x"d29c0b80",
   842 => x"f52d80d2",
   843 => x"a80b80f5",
   844 => x"2d71842b",
   845 => x"71852b07",
   846 => x"80d2b40b",
   847 => x"80f52d70",
   848 => x"822b7207",
   849 => x"80d0880c",
   850 => x"53555754",
   851 => x"9aea0480",
   852 => x"d0f40b80",
   853 => x"f52d80d1",
   854 => x"800b80f5",
   855 => x"2d71842b",
   856 => x"71852b07",
   857 => x"80d0880c",
   858 => x"545680d3",
   859 => x"c8087081",
   860 => x"06545472",
   861 => x"802e8b38",
   862 => x"80d08808",
   863 => x"810780d0",
   864 => x"880c7381",
   865 => x"2a708106",
   866 => x"51537280",
   867 => x"2e8b3880",
   868 => x"d0880882",
   869 => x"0780d088",
   870 => x"0c73822a",
   871 => x"70810651",
   872 => x"5372802e",
   873 => x"8c3880d0",
   874 => x"88088180",
   875 => x"0780d088",
   876 => x"0c80d088",
   877 => x"08fc0c86",
   878 => x"53748338",
   879 => x"845372ec",
   880 => x"0c9a8804",
   881 => x"800b80d5",
   882 => x"b40c0298",
   883 => x"050d0471",
   884 => x"980c04ff",
   885 => x"b00880d5",
   886 => x"b40c0481",
   887 => x"0bffb00c",
   888 => x"04800bff",
   889 => x"b00c0402",
   890 => x"f4050d9c",
   891 => x"f50480d5",
   892 => x"b40881f0",
   893 => x"2e098106",
   894 => x"8a38810b",
   895 => x"80d3c00c",
   896 => x"9cf50480",
   897 => x"d5b40881",
   898 => x"e02e0981",
   899 => x"068a3881",
   900 => x"0b80d3c4",
   901 => x"0c9cf504",
   902 => x"80d5b408",
   903 => x"5280d3c4",
   904 => x"08802e89",
   905 => x"3880d5b4",
   906 => x"08818005",
   907 => x"5271842c",
   908 => x"728f0653",
   909 => x"5380d3c0",
   910 => x"08802e9a",
   911 => x"38728429",
   912 => x"80d38005",
   913 => x"72138171",
   914 => x"2b700973",
   915 => x"0806730c",
   916 => x"5153539c",
   917 => x"e9047284",
   918 => x"2980d380",
   919 => x"05721383",
   920 => x"712b7208",
   921 => x"07720c53",
   922 => x"53800b80",
   923 => x"d3c40c80",
   924 => x"0b80d3c0",
   925 => x"0c80d5dc",
   926 => x"519dfc2d",
   927 => x"80d5b408",
   928 => x"ff24feea",
   929 => x"38800b80",
   930 => x"d5b40c02",
   931 => x"8c050d04",
   932 => x"02f8050d",
   933 => x"80d38052",
   934 => x"8f518072",
   935 => x"70840554",
   936 => x"0cff1151",
   937 => x"708025f2",
   938 => x"38028805",
   939 => x"0d0402f0",
   940 => x"050d7551",
   941 => x"9be12d70",
   942 => x"822cfc06",
   943 => x"80d38011",
   944 => x"72109e06",
   945 => x"71087072",
   946 => x"2a708306",
   947 => x"82742b70",
   948 => x"09740676",
   949 => x"0c545156",
   950 => x"57535153",
   951 => x"9bdb2d71",
   952 => x"80d5b40c",
   953 => x"0290050d",
   954 => x"0402fc05",
   955 => x"0d725180",
   956 => x"710c800b",
   957 => x"84120c02",
   958 => x"84050d04",
   959 => x"02f0050d",
   960 => x"75700884",
   961 => x"12085353",
   962 => x"53ff5471",
   963 => x"712ea838",
   964 => x"9be12d84",
   965 => x"13087084",
   966 => x"29148811",
   967 => x"70087081",
   968 => x"ff068418",
   969 => x"08811187",
   970 => x"06841a0c",
   971 => x"53515551",
   972 => x"51519bdb",
   973 => x"2d715473",
   974 => x"80d5b40c",
   975 => x"0290050d",
   976 => x"0402f405",
   977 => x"0d9be12d",
   978 => x"e008708b",
   979 => x"2a708106",
   980 => x"51525370",
   981 => x"802ea138",
   982 => x"80d5dc08",
   983 => x"70842980",
   984 => x"d5e40574",
   985 => x"81ff0671",
   986 => x"0c515180",
   987 => x"d5dc0881",
   988 => x"11870680",
   989 => x"d5dc0c51",
   990 => x"728c2c83",
   991 => x"ff0680d6",
   992 => x"840c800b",
   993 => x"80d6880c",
   994 => x"9bd32d9b",
   995 => x"db2d028c",
   996 => x"050d0402",
   997 => x"fc050d9b",
   998 => x"e12d810b",
   999 => x"80d6880c",
  1000 => x"9bdb2d80",
  1001 => x"d6880851",
  1002 => x"70f93802",
  1003 => x"84050d04",
  1004 => x"02fc050d",
  1005 => x"80d5dc51",
  1006 => x"9de92d9d",
  1007 => x"902d9ec1",
  1008 => x"519bcf2d",
  1009 => x"0284050d",
  1010 => x"0402fc05",
  1011 => x"0d8fcf51",
  1012 => x"86ec2dff",
  1013 => x"11517080",
  1014 => x"25f63802",
  1015 => x"84050d04",
  1016 => x"80d69008",
  1017 => x"80d5b40c",
  1018 => x"0402fc05",
  1019 => x"0d810b80",
  1020 => x"d3f40c81",
  1021 => x"51858d2d",
  1022 => x"0284050d",
  1023 => x"0402fc05",
  1024 => x"0da08704",
  1025 => x"9be72d80",
  1026 => x"f6519dae",
  1027 => x"2d80d5b4",
  1028 => x"08f23880",
  1029 => x"da519dae",
  1030 => x"2d80d5b4",
  1031 => x"08e63880",
  1032 => x"d3f00851",
  1033 => x"9dae2d80",
  1034 => x"d5b408d8",
  1035 => x"3880d5b4",
  1036 => x"0880d3f4",
  1037 => x"0c80d5b4",
  1038 => x"0851858d",
  1039 => x"2d028405",
  1040 => x"0d0402ec",
  1041 => x"050d7654",
  1042 => x"8052870b",
  1043 => x"881580f5",
  1044 => x"2d565374",
  1045 => x"72248338",
  1046 => x"a0537251",
  1047 => x"83842d81",
  1048 => x"128b1580",
  1049 => x"f52d5452",
  1050 => x"727225de",
  1051 => x"38029405",
  1052 => x"0d0402f0",
  1053 => x"050d80d6",
  1054 => x"90085481",
  1055 => x"f92d800b",
  1056 => x"80d6940c",
  1057 => x"7308802e",
  1058 => x"81893882",
  1059 => x"0b80d5c8",
  1060 => x"0c80d694",
  1061 => x"088f0680",
  1062 => x"d5c40c73",
  1063 => x"08527183",
  1064 => x"2e963871",
  1065 => x"83268938",
  1066 => x"71812eb0",
  1067 => x"38a1fc04",
  1068 => x"71852ea0",
  1069 => x"38a1fc04",
  1070 => x"881480f5",
  1071 => x"2d841508",
  1072 => x"80cecc53",
  1073 => x"545286c5",
  1074 => x"2d718429",
  1075 => x"13700852",
  1076 => x"52a28004",
  1077 => x"7351a0c2",
  1078 => x"2da1fc04",
  1079 => x"80d3c808",
  1080 => x"8815082c",
  1081 => x"70810651",
  1082 => x"5271802e",
  1083 => x"883880ce",
  1084 => x"d051a1f9",
  1085 => x"0480ced4",
  1086 => x"5186c52d",
  1087 => x"84140851",
  1088 => x"86c52d80",
  1089 => x"d6940881",
  1090 => x"0580d694",
  1091 => x"0c8c1454",
  1092 => x"a1840402",
  1093 => x"90050d04",
  1094 => x"7180d690",
  1095 => x"0ca0f22d",
  1096 => x"80d69408",
  1097 => x"ff0580d6",
  1098 => x"980c0402",
  1099 => x"e8050d80",
  1100 => x"d6900880",
  1101 => x"d69c0857",
  1102 => x"5580f651",
  1103 => x"9dae2d80",
  1104 => x"d5b40881",
  1105 => x"2a708106",
  1106 => x"51527180",
  1107 => x"2ea238a2",
  1108 => x"d5049be7",
  1109 => x"2d80f651",
  1110 => x"9dae2d80",
  1111 => x"d5b408f2",
  1112 => x"3880d3f4",
  1113 => x"08813270",
  1114 => x"80d3f40c",
  1115 => x"51858d2d",
  1116 => x"800b80d6",
  1117 => x"8c0c8c51",
  1118 => x"9dae2d80",
  1119 => x"d5b40881",
  1120 => x"2a708106",
  1121 => x"51527180",
  1122 => x"2e80d138",
  1123 => x"80d3cc08",
  1124 => x"80d3e008",
  1125 => x"80d3cc0c",
  1126 => x"80d3e00c",
  1127 => x"80d3d008",
  1128 => x"80d3e408",
  1129 => x"80d3d00c",
  1130 => x"80d3e40c",
  1131 => x"80d3d408",
  1132 => x"80d3e808",
  1133 => x"80d3d40c",
  1134 => x"80d3e80c",
  1135 => x"80d3d808",
  1136 => x"80d3ec08",
  1137 => x"80d3d80c",
  1138 => x"80d3ec0c",
  1139 => x"80d3dc08",
  1140 => x"80d3f008",
  1141 => x"80d3dc0c",
  1142 => x"80d3f00c",
  1143 => x"80d68408",
  1144 => x"a0065280",
  1145 => x"72259638",
  1146 => x"9fc92d9b",
  1147 => x"e72d80d3",
  1148 => x"f4088132",
  1149 => x"7080d3f4",
  1150 => x"0c51858d",
  1151 => x"2d80d3f4",
  1152 => x"0882ef38",
  1153 => x"80d3e008",
  1154 => x"519dae2d",
  1155 => x"80d5b408",
  1156 => x"802e8b38",
  1157 => x"80d68c08",
  1158 => x"810780d6",
  1159 => x"8c0c80d3",
  1160 => x"e408519d",
  1161 => x"ae2d80d5",
  1162 => x"b408802e",
  1163 => x"8b3880d6",
  1164 => x"8c088207",
  1165 => x"80d68c0c",
  1166 => x"80d3e808",
  1167 => x"519dae2d",
  1168 => x"80d5b408",
  1169 => x"802e8b38",
  1170 => x"80d68c08",
  1171 => x"840780d6",
  1172 => x"8c0c80d3",
  1173 => x"ec08519d",
  1174 => x"ae2d80d5",
  1175 => x"b408802e",
  1176 => x"8b3880d6",
  1177 => x"8c088807",
  1178 => x"80d68c0c",
  1179 => x"80d3f008",
  1180 => x"519dae2d",
  1181 => x"80d5b408",
  1182 => x"802e8b38",
  1183 => x"80d68c08",
  1184 => x"900780d6",
  1185 => x"8c0c80d3",
  1186 => x"cc08519d",
  1187 => x"ae2d80d5",
  1188 => x"b408802e",
  1189 => x"8c3880d6",
  1190 => x"8c088280",
  1191 => x"0780d68c",
  1192 => x"0c80d3d0",
  1193 => x"08519dae",
  1194 => x"2d80d5b4",
  1195 => x"08802e8c",
  1196 => x"3880d68c",
  1197 => x"08848007",
  1198 => x"80d68c0c",
  1199 => x"80d3d408",
  1200 => x"519dae2d",
  1201 => x"80d5b408",
  1202 => x"802e8c38",
  1203 => x"80d68c08",
  1204 => x"88800780",
  1205 => x"d68c0c80",
  1206 => x"d3d80851",
  1207 => x"9dae2d80",
  1208 => x"d5b40880",
  1209 => x"2e8c3880",
  1210 => x"d68c0890",
  1211 => x"800780d6",
  1212 => x"8c0c80d3",
  1213 => x"dc08519d",
  1214 => x"ae2d80d5",
  1215 => x"b408802e",
  1216 => x"8c3880d6",
  1217 => x"8c08a080",
  1218 => x"0780d68c",
  1219 => x"0c94519d",
  1220 => x"ae2d80d5",
  1221 => x"b4085291",
  1222 => x"519dae2d",
  1223 => x"7180d5b4",
  1224 => x"08065280",
  1225 => x"e6519dae",
  1226 => x"2d7180d5",
  1227 => x"b4080652",
  1228 => x"71802e8d",
  1229 => x"3880d68c",
  1230 => x"08848080",
  1231 => x"0780d68c",
  1232 => x"0c80fe51",
  1233 => x"9dae2d80",
  1234 => x"d5b40852",
  1235 => x"87519dae",
  1236 => x"2d7180d5",
  1237 => x"b4080752",
  1238 => x"71802e8d",
  1239 => x"3880d68c",
  1240 => x"08888080",
  1241 => x"0780d68c",
  1242 => x"0c80d68c",
  1243 => x"08ed0cae",
  1244 => x"fd049451",
  1245 => x"9dae2d80",
  1246 => x"d5b40852",
  1247 => x"91519dae",
  1248 => x"2d7180d5",
  1249 => x"b4080652",
  1250 => x"80e6519d",
  1251 => x"ae2d7180",
  1252 => x"d5b40806",
  1253 => x"5271802e",
  1254 => x"8d3880d6",
  1255 => x"8c088480",
  1256 => x"800780d6",
  1257 => x"8c0c80fe",
  1258 => x"519dae2d",
  1259 => x"80d5b408",
  1260 => x"5287519d",
  1261 => x"ae2d7180",
  1262 => x"d5b40807",
  1263 => x"5271802e",
  1264 => x"8d3880d6",
  1265 => x"8c088880",
  1266 => x"800780d6",
  1267 => x"8c0c80d6",
  1268 => x"8c08ed0c",
  1269 => x"81f5519d",
  1270 => x"ae2d80d5",
  1271 => x"b408812a",
  1272 => x"70810651",
  1273 => x"5271a438",
  1274 => x"80d3e008",
  1275 => x"519dae2d",
  1276 => x"80d5b408",
  1277 => x"812a7081",
  1278 => x"06515271",
  1279 => x"8e3880d6",
  1280 => x"84088106",
  1281 => x"52807225",
  1282 => x"80c23880",
  1283 => x"d6840881",
  1284 => x"06528072",
  1285 => x"2584389f",
  1286 => x"c92d80d6",
  1287 => x"98085271",
  1288 => x"802e8a38",
  1289 => x"ff1280d6",
  1290 => x"980ca8cc",
  1291 => x"0480d694",
  1292 => x"081080d6",
  1293 => x"94080570",
  1294 => x"84291651",
  1295 => x"52881208",
  1296 => x"802e8938",
  1297 => x"ff518812",
  1298 => x"0852712d",
  1299 => x"81f2519d",
  1300 => x"ae2d80d5",
  1301 => x"b408812a",
  1302 => x"70810651",
  1303 => x"5271a438",
  1304 => x"80d3e408",
  1305 => x"519dae2d",
  1306 => x"80d5b408",
  1307 => x"812a7081",
  1308 => x"06515271",
  1309 => x"8e3880d6",
  1310 => x"84088206",
  1311 => x"52807225",
  1312 => x"80c33880",
  1313 => x"d6840882",
  1314 => x"06528072",
  1315 => x"2584389f",
  1316 => x"c92d80d6",
  1317 => x"9408ff11",
  1318 => x"80d69808",
  1319 => x"56535373",
  1320 => x"72258a38",
  1321 => x"811480d6",
  1322 => x"980ca9c5",
  1323 => x"04721013",
  1324 => x"70842916",
  1325 => x"51528812",
  1326 => x"08802e89",
  1327 => x"38fe5188",
  1328 => x"12085271",
  1329 => x"2d81fd51",
  1330 => x"9dae2d80",
  1331 => x"d5b40881",
  1332 => x"2a708106",
  1333 => x"515271a4",
  1334 => x"3880d3e8",
  1335 => x"08519dae",
  1336 => x"2d80d5b4",
  1337 => x"08812a70",
  1338 => x"81065152",
  1339 => x"718e3880",
  1340 => x"d6840884",
  1341 => x"06528072",
  1342 => x"2580c038",
  1343 => x"80d68408",
  1344 => x"84065280",
  1345 => x"72258438",
  1346 => x"9fc92d80",
  1347 => x"d6980880",
  1348 => x"2e8a3880",
  1349 => x"0b80d698",
  1350 => x"0caabb04",
  1351 => x"80d69408",
  1352 => x"1080d694",
  1353 => x"08057084",
  1354 => x"29165152",
  1355 => x"88120880",
  1356 => x"2e8938fd",
  1357 => x"51881208",
  1358 => x"52712d81",
  1359 => x"fa519dae",
  1360 => x"2d80d5b4",
  1361 => x"08812a70",
  1362 => x"81065152",
  1363 => x"71a43880",
  1364 => x"d3ec0851",
  1365 => x"9dae2d80",
  1366 => x"d5b40881",
  1367 => x"2a708106",
  1368 => x"5152718e",
  1369 => x"3880d684",
  1370 => x"08880652",
  1371 => x"80722580",
  1372 => x"c03880d6",
  1373 => x"84088806",
  1374 => x"52807225",
  1375 => x"84389fc9",
  1376 => x"2d80d694",
  1377 => x"08ff1154",
  1378 => x"5280d698",
  1379 => x"08732589",
  1380 => x"387280d6",
  1381 => x"980cabb1",
  1382 => x"04711012",
  1383 => x"70842916",
  1384 => x"51528812",
  1385 => x"08802e89",
  1386 => x"38fc5188",
  1387 => x"12085271",
  1388 => x"2d80d698",
  1389 => x"08705354",
  1390 => x"73802e8a",
  1391 => x"388c15ff",
  1392 => x"155555ab",
  1393 => x"b804820b",
  1394 => x"80d5c80c",
  1395 => x"718f0680",
  1396 => x"d5c40c81",
  1397 => x"eb519dae",
  1398 => x"2d80d5b4",
  1399 => x"08812a70",
  1400 => x"81065152",
  1401 => x"71802ead",
  1402 => x"38740885",
  1403 => x"2e098106",
  1404 => x"a4388815",
  1405 => x"80f52dff",
  1406 => x"05527188",
  1407 => x"1681b72d",
  1408 => x"71982b52",
  1409 => x"71802588",
  1410 => x"38800b88",
  1411 => x"1681b72d",
  1412 => x"7451a0c2",
  1413 => x"2d81f451",
  1414 => x"9dae2d80",
  1415 => x"d5b40881",
  1416 => x"2a708106",
  1417 => x"51527180",
  1418 => x"2eb33874",
  1419 => x"08852e09",
  1420 => x"8106aa38",
  1421 => x"881580f5",
  1422 => x"2d810552",
  1423 => x"71881681",
  1424 => x"b72d7181",
  1425 => x"ff068b16",
  1426 => x"80f52d54",
  1427 => x"52727227",
  1428 => x"87387288",
  1429 => x"1681b72d",
  1430 => x"7451a0c2",
  1431 => x"2d80da51",
  1432 => x"9dae2d80",
  1433 => x"d5b40881",
  1434 => x"2a708106",
  1435 => x"5152718e",
  1436 => x"3880d684",
  1437 => x"08900652",
  1438 => x"80722581",
  1439 => x"bc3880d6",
  1440 => x"900880d6",
  1441 => x"84089006",
  1442 => x"53538072",
  1443 => x"2584389f",
  1444 => x"c92d80d6",
  1445 => x"98085473",
  1446 => x"802e8a38",
  1447 => x"8c13ff15",
  1448 => x"5553ad97",
  1449 => x"04720852",
  1450 => x"71822ea6",
  1451 => x"38718226",
  1452 => x"89387181",
  1453 => x"2eaa38ae",
  1454 => x"b9047183",
  1455 => x"2eb43871",
  1456 => x"842e0981",
  1457 => x"0680f238",
  1458 => x"88130851",
  1459 => x"a2982dae",
  1460 => x"b90480d6",
  1461 => x"98085188",
  1462 => x"13085271",
  1463 => x"2daeb904",
  1464 => x"810b8814",
  1465 => x"082b80d3",
  1466 => x"c8083280",
  1467 => x"d3c80cae",
  1468 => x"8d048813",
  1469 => x"80f52d81",
  1470 => x"058b1480",
  1471 => x"f52d5354",
  1472 => x"71742483",
  1473 => x"38805473",
  1474 => x"881481b7",
  1475 => x"2da0f22d",
  1476 => x"aeb90475",
  1477 => x"08802ea4",
  1478 => x"38750851",
  1479 => x"9dae2d80",
  1480 => x"d5b40881",
  1481 => x"06527180",
  1482 => x"2e8c3880",
  1483 => x"d6980851",
  1484 => x"84160852",
  1485 => x"712d8816",
  1486 => x"5675d838",
  1487 => x"8054800b",
  1488 => x"80d5c80c",
  1489 => x"738f0680",
  1490 => x"d5c40ca0",
  1491 => x"527380d6",
  1492 => x"98082e09",
  1493 => x"81069938",
  1494 => x"80d69408",
  1495 => x"ff057432",
  1496 => x"70098105",
  1497 => x"7072079f",
  1498 => x"2a917131",
  1499 => x"51515353",
  1500 => x"71518384",
  1501 => x"2d811454",
  1502 => x"8e7425c2",
  1503 => x"3880d3f4",
  1504 => x"0880d5b4",
  1505 => x"0c029805",
  1506 => x"0d0402f4",
  1507 => x"050dd452",
  1508 => x"81ff720c",
  1509 => x"71085381",
  1510 => x"ff720c72",
  1511 => x"882b83fe",
  1512 => x"80067208",
  1513 => x"7081ff06",
  1514 => x"51525381",
  1515 => x"ff720c72",
  1516 => x"7107882b",
  1517 => x"72087081",
  1518 => x"ff065152",
  1519 => x"5381ff72",
  1520 => x"0c727107",
  1521 => x"882b7208",
  1522 => x"7081ff06",
  1523 => x"720780d5",
  1524 => x"b40c5253",
  1525 => x"028c050d",
  1526 => x"0402f405",
  1527 => x"0d747671",
  1528 => x"81ff06d4",
  1529 => x"0c535380",
  1530 => x"d6a00885",
  1531 => x"3871892b",
  1532 => x"5271982a",
  1533 => x"d40c7190",
  1534 => x"2a7081ff",
  1535 => x"06d40c51",
  1536 => x"71882a70",
  1537 => x"81ff06d4",
  1538 => x"0c517181",
  1539 => x"ff06d40c",
  1540 => x"72902a70",
  1541 => x"81ff06d4",
  1542 => x"0c51d408",
  1543 => x"7081ff06",
  1544 => x"515182b8",
  1545 => x"bf527081",
  1546 => x"ff2e0981",
  1547 => x"06943881",
  1548 => x"ff0bd40c",
  1549 => x"d4087081",
  1550 => x"ff06ff14",
  1551 => x"54515171",
  1552 => x"e5387080",
  1553 => x"d5b40c02",
  1554 => x"8c050d04",
  1555 => x"02fc050d",
  1556 => x"81c75181",
  1557 => x"ff0bd40c",
  1558 => x"ff115170",
  1559 => x"8025f438",
  1560 => x"0284050d",
  1561 => x"0402f405",
  1562 => x"0d81ff0b",
  1563 => x"d40c9353",
  1564 => x"805287fc",
  1565 => x"80c151af",
  1566 => x"d92d80d5",
  1567 => x"b4088b38",
  1568 => x"81ff0bd4",
  1569 => x"0c8153b1",
  1570 => x"9304b0cc",
  1571 => x"2dff1353",
  1572 => x"72de3872",
  1573 => x"80d5b40c",
  1574 => x"028c050d",
  1575 => x"0402ec05",
  1576 => x"0d810b80",
  1577 => x"d6a00c84",
  1578 => x"54d00870",
  1579 => x"8f2a7081",
  1580 => x"06515153",
  1581 => x"72f33872",
  1582 => x"d00cb0cc",
  1583 => x"2d80ced8",
  1584 => x"5186c52d",
  1585 => x"d008708f",
  1586 => x"2a708106",
  1587 => x"51515372",
  1588 => x"f338810b",
  1589 => x"d00cb153",
  1590 => x"805284d4",
  1591 => x"80c051af",
  1592 => x"d92d80d5",
  1593 => x"b408812e",
  1594 => x"93387282",
  1595 => x"2ebf38ff",
  1596 => x"135372e4",
  1597 => x"38ff1454",
  1598 => x"73ffae38",
  1599 => x"b0cc2d83",
  1600 => x"aa52849c",
  1601 => x"80c851af",
  1602 => x"d92d80d5",
  1603 => x"b408812e",
  1604 => x"09810693",
  1605 => x"38af8a2d",
  1606 => x"80d5b408",
  1607 => x"83ffff06",
  1608 => x"537283aa",
  1609 => x"2e9f38b0",
  1610 => x"e52db2c0",
  1611 => x"0480cee4",
  1612 => x"5186c52d",
  1613 => x"8053b495",
  1614 => x"0480cefc",
  1615 => x"5186c52d",
  1616 => x"8054b3e6",
  1617 => x"0481ff0b",
  1618 => x"d40cb154",
  1619 => x"b0cc2d8f",
  1620 => x"cf538052",
  1621 => x"87fc80f7",
  1622 => x"51afd92d",
  1623 => x"80d5b408",
  1624 => x"5580d5b4",
  1625 => x"08812e09",
  1626 => x"81069c38",
  1627 => x"81ff0bd4",
  1628 => x"0c820a52",
  1629 => x"849c80e9",
  1630 => x"51afd92d",
  1631 => x"80d5b408",
  1632 => x"802e8d38",
  1633 => x"b0cc2dff",
  1634 => x"135372c6",
  1635 => x"38b3d904",
  1636 => x"81ff0bd4",
  1637 => x"0c80d5b4",
  1638 => x"085287fc",
  1639 => x"80fa51af",
  1640 => x"d92d80d5",
  1641 => x"b408b238",
  1642 => x"81ff0bd4",
  1643 => x"0cd40853",
  1644 => x"81ff0bd4",
  1645 => x"0c81ff0b",
  1646 => x"d40c81ff",
  1647 => x"0bd40c81",
  1648 => x"ff0bd40c",
  1649 => x"72862a70",
  1650 => x"81067656",
  1651 => x"51537296",
  1652 => x"3880d5b4",
  1653 => x"0854b3e6",
  1654 => x"0473822e",
  1655 => x"fedb38ff",
  1656 => x"145473fe",
  1657 => x"e7387380",
  1658 => x"d6a00c73",
  1659 => x"8b388152",
  1660 => x"87fc80d0",
  1661 => x"51afd92d",
  1662 => x"81ff0bd4",
  1663 => x"0cd00870",
  1664 => x"8f2a7081",
  1665 => x"06515153",
  1666 => x"72f33872",
  1667 => x"d00c81ff",
  1668 => x"0bd40c81",
  1669 => x"537280d5",
  1670 => x"b40c0294",
  1671 => x"050d0402",
  1672 => x"e8050d78",
  1673 => x"55805681",
  1674 => x"ff0bd40c",
  1675 => x"d008708f",
  1676 => x"2a708106",
  1677 => x"51515372",
  1678 => x"f3388281",
  1679 => x"0bd00c81",
  1680 => x"ff0bd40c",
  1681 => x"775287fc",
  1682 => x"80d151af",
  1683 => x"d92d80db",
  1684 => x"c6df5480",
  1685 => x"d5b40880",
  1686 => x"2e8b3880",
  1687 => x"cf9c5186",
  1688 => x"c52db5b9",
  1689 => x"0481ff0b",
  1690 => x"d40cd408",
  1691 => x"7081ff06",
  1692 => x"51537281",
  1693 => x"fe2e0981",
  1694 => x"069e3880",
  1695 => x"ff53af8a",
  1696 => x"2d80d5b4",
  1697 => x"08757084",
  1698 => x"05570cff",
  1699 => x"13537280",
  1700 => x"25ec3881",
  1701 => x"56b59e04",
  1702 => x"ff145473",
  1703 => x"c83881ff",
  1704 => x"0bd40c81",
  1705 => x"ff0bd40c",
  1706 => x"d008708f",
  1707 => x"2a708106",
  1708 => x"51515372",
  1709 => x"f33872d0",
  1710 => x"0c7580d5",
  1711 => x"b40c0298",
  1712 => x"050d0402",
  1713 => x"e8050d77",
  1714 => x"797b5855",
  1715 => x"55805372",
  1716 => x"7625a338",
  1717 => x"74708105",
  1718 => x"5680f52d",
  1719 => x"74708105",
  1720 => x"5680f52d",
  1721 => x"52527171",
  1722 => x"2e863881",
  1723 => x"51b5f804",
  1724 => x"811353b5",
  1725 => x"cf048051",
  1726 => x"7080d5b4",
  1727 => x"0c029805",
  1728 => x"0d0402ec",
  1729 => x"050d7655",
  1730 => x"74802e80",
  1731 => x"c4389a15",
  1732 => x"80e02d51",
  1733 => x"80c4a22d",
  1734 => x"80d5b408",
  1735 => x"80d5b408",
  1736 => x"80dcd40c",
  1737 => x"80d5b408",
  1738 => x"545480dc",
  1739 => x"b008802e",
  1740 => x"9b389415",
  1741 => x"80e02d51",
  1742 => x"80c4a22d",
  1743 => x"80d5b408",
  1744 => x"902b83ff",
  1745 => x"f00a0670",
  1746 => x"75075153",
  1747 => x"7280dcd4",
  1748 => x"0c80dcd4",
  1749 => x"08537280",
  1750 => x"2e9d3880",
  1751 => x"dca808fe",
  1752 => x"14712980",
  1753 => x"dcbc0805",
  1754 => x"80dcd80c",
  1755 => x"70842b80",
  1756 => x"dcb40c54",
  1757 => x"b7a50480",
  1758 => x"dcc00880",
  1759 => x"dcd40c80",
  1760 => x"dcc40880",
  1761 => x"dcd80c80",
  1762 => x"dcb00880",
  1763 => x"2e8b3880",
  1764 => x"dca80884",
  1765 => x"2b53b7a0",
  1766 => x"0480dcc8",
  1767 => x"08842b53",
  1768 => x"7280dcb4",
  1769 => x"0c029405",
  1770 => x"0d0402d8",
  1771 => x"050d800b",
  1772 => x"80dcb00c",
  1773 => x"8454b19d",
  1774 => x"2d80d5b4",
  1775 => x"08802e97",
  1776 => x"3880d6a4",
  1777 => x"528051b4",
  1778 => x"9f2d80d5",
  1779 => x"b408802e",
  1780 => x"8638fe54",
  1781 => x"b7df04ff",
  1782 => x"14547380",
  1783 => x"24d83873",
  1784 => x"8d3880cf",
  1785 => x"ac5186c5",
  1786 => x"2d7355bd",
  1787 => x"b5048056",
  1788 => x"810b80dc",
  1789 => x"dc0c8853",
  1790 => x"80cfc052",
  1791 => x"80d6da51",
  1792 => x"b5c32d80",
  1793 => x"d5b40876",
  1794 => x"2e098106",
  1795 => x"893880d5",
  1796 => x"b40880dc",
  1797 => x"dc0c8853",
  1798 => x"80cfcc52",
  1799 => x"80d6f651",
  1800 => x"b5c32d80",
  1801 => x"d5b40889",
  1802 => x"3880d5b4",
  1803 => x"0880dcdc",
  1804 => x"0c80dcdc",
  1805 => x"08802e81",
  1806 => x"823880d9",
  1807 => x"ea0b80f5",
  1808 => x"2d80d9eb",
  1809 => x"0b80f52d",
  1810 => x"71982b71",
  1811 => x"902b0780",
  1812 => x"d9ec0b80",
  1813 => x"f52d7088",
  1814 => x"2b720780",
  1815 => x"d9ed0b80",
  1816 => x"f52d7107",
  1817 => x"80daa20b",
  1818 => x"80f52d80",
  1819 => x"daa30b80",
  1820 => x"f52d7188",
  1821 => x"2b07535f",
  1822 => x"54525a56",
  1823 => x"57557381",
  1824 => x"abaa2e09",
  1825 => x"81068f38",
  1826 => x"755180c3",
  1827 => x"f12d80d5",
  1828 => x"b40856b9",
  1829 => x"a4047382",
  1830 => x"d4d52e88",
  1831 => x"3880cfd8",
  1832 => x"51b9f004",
  1833 => x"80d6a452",
  1834 => x"7551b49f",
  1835 => x"2d80d5b4",
  1836 => x"085580d5",
  1837 => x"b408802e",
  1838 => x"83fb3888",
  1839 => x"5380cfcc",
  1840 => x"5280d6f6",
  1841 => x"51b5c32d",
  1842 => x"80d5b408",
  1843 => x"8a38810b",
  1844 => x"80dcb00c",
  1845 => x"b9f60488",
  1846 => x"5380cfc0",
  1847 => x"5280d6da",
  1848 => x"51b5c32d",
  1849 => x"80d5b408",
  1850 => x"802e8b38",
  1851 => x"80cfec51",
  1852 => x"86c52dba",
  1853 => x"d50480da",
  1854 => x"a20b80f5",
  1855 => x"2d547380",
  1856 => x"d52e0981",
  1857 => x"0680ce38",
  1858 => x"80daa30b",
  1859 => x"80f52d54",
  1860 => x"7381aa2e",
  1861 => x"098106bd",
  1862 => x"38800b80",
  1863 => x"d6a40b80",
  1864 => x"f52d5654",
  1865 => x"7481e92e",
  1866 => x"83388154",
  1867 => x"7481eb2e",
  1868 => x"8c388055",
  1869 => x"73752e09",
  1870 => x"810682f9",
  1871 => x"3880d6af",
  1872 => x"0b80f52d",
  1873 => x"55748e38",
  1874 => x"80d6b00b",
  1875 => x"80f52d54",
  1876 => x"73822e86",
  1877 => x"388055bd",
  1878 => x"b50480d6",
  1879 => x"b10b80f5",
  1880 => x"2d7080dc",
  1881 => x"a80cff05",
  1882 => x"80dcac0c",
  1883 => x"80d6b20b",
  1884 => x"80f52d80",
  1885 => x"d6b30b80",
  1886 => x"f52d5876",
  1887 => x"05778280",
  1888 => x"29057080",
  1889 => x"dcb80c80",
  1890 => x"d6b40b80",
  1891 => x"f52d7080",
  1892 => x"dccc0c80",
  1893 => x"dcb00859",
  1894 => x"57587680",
  1895 => x"2e81b738",
  1896 => x"885380cf",
  1897 => x"cc5280d6",
  1898 => x"f651b5c3",
  1899 => x"2d80d5b4",
  1900 => x"08828238",
  1901 => x"80dca808",
  1902 => x"70842b80",
  1903 => x"dcb40c70",
  1904 => x"80dcc80c",
  1905 => x"80d6c90b",
  1906 => x"80f52d80",
  1907 => x"d6c80b80",
  1908 => x"f52d7182",
  1909 => x"80290580",
  1910 => x"d6ca0b80",
  1911 => x"f52d7084",
  1912 => x"80802912",
  1913 => x"80d6cb0b",
  1914 => x"80f52d70",
  1915 => x"81800a29",
  1916 => x"127080dc",
  1917 => x"d00c80dc",
  1918 => x"cc087129",
  1919 => x"80dcb808",
  1920 => x"057080dc",
  1921 => x"bc0c80d6",
  1922 => x"d10b80f5",
  1923 => x"2d80d6d0",
  1924 => x"0b80f52d",
  1925 => x"71828029",
  1926 => x"0580d6d2",
  1927 => x"0b80f52d",
  1928 => x"70848080",
  1929 => x"291280d6",
  1930 => x"d30b80f5",
  1931 => x"2d70982b",
  1932 => x"81f00a06",
  1933 => x"72057080",
  1934 => x"dcc00cfe",
  1935 => x"117e2977",
  1936 => x"0580dcc4",
  1937 => x"0c525952",
  1938 => x"43545e51",
  1939 => x"5259525d",
  1940 => x"575957bd",
  1941 => x"ae0480d6",
  1942 => x"b60b80f5",
  1943 => x"2d80d6b5",
  1944 => x"0b80f52d",
  1945 => x"71828029",
  1946 => x"057080dc",
  1947 => x"b40c70a0",
  1948 => x"2983ff05",
  1949 => x"70892a70",
  1950 => x"80dcc80c",
  1951 => x"80d6bb0b",
  1952 => x"80f52d80",
  1953 => x"d6ba0b80",
  1954 => x"f52d7182",
  1955 => x"80290570",
  1956 => x"80dcd00c",
  1957 => x"7b71291e",
  1958 => x"7080dcc4",
  1959 => x"0c7d80dc",
  1960 => x"c00c7305",
  1961 => x"80dcbc0c",
  1962 => x"555e5151",
  1963 => x"55558051",
  1964 => x"b6822d81",
  1965 => x"557480d5",
  1966 => x"b40c02a8",
  1967 => x"050d0402",
  1968 => x"ec050d76",
  1969 => x"70872c71",
  1970 => x"80ff0655",
  1971 => x"565480dc",
  1972 => x"b0088a38",
  1973 => x"73882c74",
  1974 => x"81ff0654",
  1975 => x"5580d6a4",
  1976 => x"5280dcb8",
  1977 => x"081551b4",
  1978 => x"9f2d80d5",
  1979 => x"b4085480",
  1980 => x"d5b40880",
  1981 => x"2eba3880",
  1982 => x"dcb00880",
  1983 => x"2e9b3872",
  1984 => x"842980d6",
  1985 => x"a4057008",
  1986 => x"525380c3",
  1987 => x"f12d80d5",
  1988 => x"b408f00a",
  1989 => x"0653beae",
  1990 => x"04721080",
  1991 => x"d6a40570",
  1992 => x"80e02d52",
  1993 => x"5380c4a2",
  1994 => x"2d80d5b4",
  1995 => x"08537254",
  1996 => x"7380d5b4",
  1997 => x"0c029405",
  1998 => x"0d0402e0",
  1999 => x"050d7970",
  2000 => x"842c80dc",
  2001 => x"d8080571",
  2002 => x"8f065255",
  2003 => x"53728a38",
  2004 => x"80d6a452",
  2005 => x"7351b49f",
  2006 => x"2d72a029",
  2007 => x"80d6a405",
  2008 => x"54807480",
  2009 => x"f52d5653",
  2010 => x"74732e83",
  2011 => x"38815374",
  2012 => x"81e52e81",
  2013 => x"f5388170",
  2014 => x"74065458",
  2015 => x"72802e81",
  2016 => x"e9388b14",
  2017 => x"80f52d70",
  2018 => x"832a7906",
  2019 => x"5856769c",
  2020 => x"3880d3f8",
  2021 => x"08537289",
  2022 => x"387280da",
  2023 => x"a40b81b7",
  2024 => x"2d7680d3",
  2025 => x"f80c7353",
  2026 => x"80c0ec04",
  2027 => x"758f2e09",
  2028 => x"810681b6",
  2029 => x"38749f06",
  2030 => x"8d2980da",
  2031 => x"97115153",
  2032 => x"811480f5",
  2033 => x"2d737081",
  2034 => x"055581b7",
  2035 => x"2d831480",
  2036 => x"f52d7370",
  2037 => x"81055581",
  2038 => x"b72d8514",
  2039 => x"80f52d73",
  2040 => x"70810555",
  2041 => x"81b72d87",
  2042 => x"1480f52d",
  2043 => x"73708105",
  2044 => x"5581b72d",
  2045 => x"891480f5",
  2046 => x"2d737081",
  2047 => x"055581b7",
  2048 => x"2d8e1480",
  2049 => x"f52d7370",
  2050 => x"81055581",
  2051 => x"b72d9014",
  2052 => x"80f52d73",
  2053 => x"70810555",
  2054 => x"81b72d92",
  2055 => x"1480f52d",
  2056 => x"73708105",
  2057 => x"5581b72d",
  2058 => x"941480f5",
  2059 => x"2d737081",
  2060 => x"055581b7",
  2061 => x"2d961480",
  2062 => x"f52d7370",
  2063 => x"81055581",
  2064 => x"b72d9814",
  2065 => x"80f52d73",
  2066 => x"70810555",
  2067 => x"81b72d9c",
  2068 => x"1480f52d",
  2069 => x"73708105",
  2070 => x"5581b72d",
  2071 => x"9e1480f5",
  2072 => x"2d7381b7",
  2073 => x"2d7780d3",
  2074 => x"f80c8053",
  2075 => x"7280d5b4",
  2076 => x"0c02a005",
  2077 => x"0d0402cc",
  2078 => x"050d7e60",
  2079 => x"5e5a800b",
  2080 => x"80dcd408",
  2081 => x"80dcd808",
  2082 => x"595c5680",
  2083 => x"5880dcb4",
  2084 => x"08782e81",
  2085 => x"bc38778f",
  2086 => x"06a01757",
  2087 => x"54739138",
  2088 => x"80d6a452",
  2089 => x"76518117",
  2090 => x"57b49f2d",
  2091 => x"80d6a456",
  2092 => x"807680f5",
  2093 => x"2d565474",
  2094 => x"742e8338",
  2095 => x"81547481",
  2096 => x"e52e8181",
  2097 => x"38817075",
  2098 => x"06555c73",
  2099 => x"802e80f5",
  2100 => x"388b1680",
  2101 => x"f52d9806",
  2102 => x"597880e9",
  2103 => x"388b537c",
  2104 => x"527551b5",
  2105 => x"c32d80d5",
  2106 => x"b40880d9",
  2107 => x"389c1608",
  2108 => x"5180c3f1",
  2109 => x"2d80d5b4",
  2110 => x"08841b0c",
  2111 => x"9a1680e0",
  2112 => x"2d5180c4",
  2113 => x"a22d80d5",
  2114 => x"b40880d5",
  2115 => x"b408881c",
  2116 => x"0c80d5b4",
  2117 => x"08555580",
  2118 => x"dcb00880",
  2119 => x"2e9a3894",
  2120 => x"1680e02d",
  2121 => x"5180c4a2",
  2122 => x"2d80d5b4",
  2123 => x"08902b83",
  2124 => x"fff00a06",
  2125 => x"70165154",
  2126 => x"73881b0c",
  2127 => x"787a0c7b",
  2128 => x"5480c38e",
  2129 => x"04811858",
  2130 => x"80dcb408",
  2131 => x"7826fec6",
  2132 => x"3880dcb0",
  2133 => x"08802eb4",
  2134 => x"387a51bd",
  2135 => x"bf2d80d5",
  2136 => x"b40880d5",
  2137 => x"b40880ff",
  2138 => x"fffff806",
  2139 => x"555b7380",
  2140 => x"fffffff8",
  2141 => x"2e963880",
  2142 => x"d5b408fe",
  2143 => x"0580dca8",
  2144 => x"082980dc",
  2145 => x"bc080557",
  2146 => x"80c18b04",
  2147 => x"80547380",
  2148 => x"d5b40c02",
  2149 => x"b4050d04",
  2150 => x"02f4050d",
  2151 => x"74700881",
  2152 => x"05710c70",
  2153 => x"0880dcac",
  2154 => x"08065353",
  2155 => x"718f3888",
  2156 => x"130851bd",
  2157 => x"bf2d80d5",
  2158 => x"b4088814",
  2159 => x"0c810b80",
  2160 => x"d5b40c02",
  2161 => x"8c050d04",
  2162 => x"02f0050d",
  2163 => x"75881108",
  2164 => x"fe0580dc",
  2165 => x"a8082980",
  2166 => x"dcbc0811",
  2167 => x"720880dc",
  2168 => x"ac080605",
  2169 => x"79555354",
  2170 => x"54b49f2d",
  2171 => x"0290050d",
  2172 => x"0402f405",
  2173 => x"0d747088",
  2174 => x"2a83fe80",
  2175 => x"06707298",
  2176 => x"2a077288",
  2177 => x"2b87fc80",
  2178 => x"80067398",
  2179 => x"2b81f00a",
  2180 => x"06717307",
  2181 => x"0780d5b4",
  2182 => x"0c565153",
  2183 => x"51028c05",
  2184 => x"0d0402f8",
  2185 => x"050d028e",
  2186 => x"0580f52d",
  2187 => x"74882b07",
  2188 => x"7083ffff",
  2189 => x"0680d5b4",
  2190 => x"0c510288",
  2191 => x"050d0402",
  2192 => x"f4050d74",
  2193 => x"76785354",
  2194 => x"52807125",
  2195 => x"97387270",
  2196 => x"81055480",
  2197 => x"f52d7270",
  2198 => x"81055481",
  2199 => x"b72dff11",
  2200 => x"5170eb38",
  2201 => x"807281b7",
  2202 => x"2d028c05",
  2203 => x"0d0402e8",
  2204 => x"050d7756",
  2205 => x"80705654",
  2206 => x"737624b6",
  2207 => x"3880dcb4",
  2208 => x"08742eae",
  2209 => x"387351be",
  2210 => x"ba2d80d5",
  2211 => x"b40880d5",
  2212 => x"b4080981",
  2213 => x"057080d5",
  2214 => x"b408079f",
  2215 => x"2a770581",
  2216 => x"17575753",
  2217 => x"53747624",
  2218 => x"893880dc",
  2219 => x"b4087426",
  2220 => x"d4387280",
  2221 => x"d5b40c02",
  2222 => x"98050d04",
  2223 => x"02ec050d",
  2224 => x"80d5b008",
  2225 => x"175180c4",
  2226 => x"ee2d80d5",
  2227 => x"b4085580",
  2228 => x"d5b40880",
  2229 => x"2ea3388b",
  2230 => x"5380d5b4",
  2231 => x"085280da",
  2232 => x"a45180c4",
  2233 => x"bf2d80dc",
  2234 => x"e0085473",
  2235 => x"802e8a38",
  2236 => x"88155280",
  2237 => x"daa45173",
  2238 => x"2d029405",
  2239 => x"0d0402dc",
  2240 => x"050d8070",
  2241 => x"5a557480",
  2242 => x"d5b00825",
  2243 => x"b43880dc",
  2244 => x"b408752e",
  2245 => x"ac387851",
  2246 => x"beba2d80",
  2247 => x"d5b40809",
  2248 => x"81057080",
  2249 => x"d5b40807",
  2250 => x"9f2a7605",
  2251 => x"811b5b56",
  2252 => x"547480d5",
  2253 => x"b0082589",
  2254 => x"3880dcb4",
  2255 => x"087926d6",
  2256 => x"38805578",
  2257 => x"80dcb408",
  2258 => x"2781e338",
  2259 => x"7851beba",
  2260 => x"2d80d5b4",
  2261 => x"08802e81",
  2262 => x"b43880d5",
  2263 => x"b4088b05",
  2264 => x"80f52d70",
  2265 => x"842a7081",
  2266 => x"06771078",
  2267 => x"842b80da",
  2268 => x"a40b80f5",
  2269 => x"2d5c5c53",
  2270 => x"51555673",
  2271 => x"802e80ce",
  2272 => x"38741682",
  2273 => x"2b80c8d2",
  2274 => x"0b80d484",
  2275 => x"120c5477",
  2276 => x"75311080",
  2277 => x"dce41155",
  2278 => x"56907470",
  2279 => x"81055681",
  2280 => x"b72da074",
  2281 => x"81b72d76",
  2282 => x"81ff0681",
  2283 => x"16585473",
  2284 => x"802e8b38",
  2285 => x"9c5380da",
  2286 => x"a45280c7",
  2287 => x"c5048b53",
  2288 => x"80d5b408",
  2289 => x"5280dce6",
  2290 => x"165180c8",
  2291 => x"83047416",
  2292 => x"822b80c5",
  2293 => x"bc0b80d4",
  2294 => x"84120c54",
  2295 => x"7681ff06",
  2296 => x"81165854",
  2297 => x"73802e8b",
  2298 => x"389c5380",
  2299 => x"daa45280",
  2300 => x"c7fa048b",
  2301 => x"5380d5b4",
  2302 => x"08527775",
  2303 => x"311080dc",
  2304 => x"e4055176",
  2305 => x"5580c4bf",
  2306 => x"2d80c8a2",
  2307 => x"04749029",
  2308 => x"75317010",
  2309 => x"80dce405",
  2310 => x"515480d5",
  2311 => x"b4087481",
  2312 => x"b72d8119",
  2313 => x"59748b24",
  2314 => x"a43880c6",
  2315 => x"c3047490",
  2316 => x"29753170",
  2317 => x"1080dce4",
  2318 => x"058c7731",
  2319 => x"57515480",
  2320 => x"7481b72d",
  2321 => x"9e14ff16",
  2322 => x"565474f3",
  2323 => x"3802a405",
  2324 => x"0d0402fc",
  2325 => x"050d80d5",
  2326 => x"b0081351",
  2327 => x"80c4ee2d",
  2328 => x"80d5b408",
  2329 => x"802e8938",
  2330 => x"80d5b408",
  2331 => x"51b6822d",
  2332 => x"800b80d5",
  2333 => x"b00c80c5",
  2334 => x"fe2da0f2",
  2335 => x"2d028405",
  2336 => x"0d0402fc",
  2337 => x"050d7251",
  2338 => x"70fd2eb2",
  2339 => x"3870fd24",
  2340 => x"8b3870fc",
  2341 => x"2e80d038",
  2342 => x"80c9f104",
  2343 => x"70fe2eb9",
  2344 => x"3870ff2e",
  2345 => x"09810680",
  2346 => x"c83880d5",
  2347 => x"b0085170",
  2348 => x"802ebe38",
  2349 => x"ff1180d5",
  2350 => x"b00c80c9",
  2351 => x"f10480d5",
  2352 => x"b008f405",
  2353 => x"7080d5b0",
  2354 => x"0c517080",
  2355 => x"25a33880",
  2356 => x"0b80d5b0",
  2357 => x"0c80c9f1",
  2358 => x"0480d5b0",
  2359 => x"08810580",
  2360 => x"d5b00c80",
  2361 => x"c9f10480",
  2362 => x"d5b0088c",
  2363 => x"0580d5b0",
  2364 => x"0c80c5fe",
  2365 => x"2da0f22d",
  2366 => x"0284050d",
  2367 => x"0402fc05",
  2368 => x"0d800b80",
  2369 => x"d5b00c80",
  2370 => x"c5fe2d9f",
  2371 => x"e02d80d5",
  2372 => x"b40880d5",
  2373 => x"a00c80d3",
  2374 => x"fc51a298",
  2375 => x"2d028405",
  2376 => x"0d0402fc",
  2377 => x"050d810b",
  2378 => x"80d0840c",
  2379 => x"725180c9",
  2380 => x"fd2d0284",
  2381 => x"050d0402",
  2382 => x"fc050d80",
  2383 => x"0b80d084",
  2384 => x"0c725180",
  2385 => x"c9fd2d02",
  2386 => x"84050d04",
  2387 => x"7180dce0",
  2388 => x"0c040000",
  2389 => x"00ffffff",
  2390 => x"ff00ffff",
  2391 => x"ffff00ff",
  2392 => x"ffffff00",
  2393 => x"4b455953",
  2394 => x"50312020",
  2395 => x"20202000",
  2396 => x"00000000",
  2397 => x"4b455953",
  2398 => x"50322020",
  2399 => x"20202000",
  2400 => x"00000000",
  2401 => x"3d3d2056",
  2402 => x"6964656f",
  2403 => x"70616320",
  2404 => x"666f7220",
  2405 => x"5a58444f",
  2406 => x"53203d3d",
  2407 => x"00000000",
  2408 => x"3d3d3d3d",
  2409 => x"3d3d3d3d",
  2410 => x"3d3d3d3d",
  2411 => x"3d3d3d3d",
  2412 => x"3d3d3d3d",
  2413 => x"3d3d3d3d",
  2414 => x"00000000",
  2415 => x"52657365",
  2416 => x"74000000",
  2417 => x"5363616e",
  2418 => x"6c696e65",
  2419 => x"73000000",
  2420 => x"53776170",
  2421 => x"206a6f79",
  2422 => x"73746963",
  2423 => x"6b730000",
  2424 => x"4a6f696e",
  2425 => x"206a6f79",
  2426 => x"73746963",
  2427 => x"6b730000",
  2428 => x"4c6f6164",
  2429 => x"20636174",
  2430 => x"72696467",
  2431 => x"6520524f",
  2432 => x"4d201000",
  2433 => x"4c6f6164",
  2434 => x"20564443",
  2435 => x"20666f6e",
  2436 => x"74201000",
  2437 => x"45786974",
  2438 => x"00000000",
  2439 => x"436f6c6f",
  2440 => x"72206d6f",
  2441 => x"64653a20",
  2442 => x"436f6c6f",
  2443 => x"72000000",
  2444 => x"436f6c6f",
  2445 => x"72206d6f",
  2446 => x"64653a20",
  2447 => x"4d6f6e6f",
  2448 => x"6368726f",
  2449 => x"6d650000",
  2450 => x"436f6c6f",
  2451 => x"72206d6f",
  2452 => x"64653a20",
  2453 => x"47726565",
  2454 => x"6e207068",
  2455 => x"6f737068",
  2456 => x"6f720000",
  2457 => x"436f6c6f",
  2458 => x"72206d6f",
  2459 => x"64653a20",
  2460 => x"416d6265",
  2461 => x"72206d6f",
  2462 => x"6e6f6368",
  2463 => x"726f6d65",
  2464 => x"00000000",
  2465 => x"4d6f6465",
  2466 => x"3a204f64",
  2467 => x"79737365",
  2468 => x"79322028",
  2469 => x"4e545343",
  2470 => x"29000000",
  2471 => x"4d6f6465",
  2472 => x"3a205669",
  2473 => x"64656f70",
  2474 => x"61632028",
  2475 => x"50414c29",
  2476 => x"00000000",
  2477 => x"3d3d2056",
  2478 => x"6964656f",
  2479 => x"70616320",
  2480 => x"666f7220",
  2481 => x"5a58554e",
  2482 => x"4f203d3d",
  2483 => x"00000000",
  2484 => x"5a58554e",
  2485 => x"4f3a2073",
  2486 => x"696e676c",
  2487 => x"65206a6f",
  2488 => x"79737469",
  2489 => x"636b0000",
  2490 => x"5a58554e",
  2491 => x"4f3a2032",
  2492 => x"206a6f79",
  2493 => x"73746963",
  2494 => x"6b207370",
  2495 => x"6c697474",
  2496 => x"65720000",
  2497 => x"5a58554e",
  2498 => x"4f3a2032",
  2499 => x"206a6f79",
  2500 => x"73746963",
  2501 => x"6b205647",
  2502 => x"41324d00",
  2503 => x"524f4d20",
  2504 => x"6c6f6164",
  2505 => x"696e6720",
  2506 => x"6661696c",
  2507 => x"65640000",
  2508 => x"4f4b0000",
  2509 => x"496e6974",
  2510 => x"69616c69",
  2511 => x"7a696e67",
  2512 => x"20534420",
  2513 => x"63617264",
  2514 => x"0a000000",
  2515 => x"16200000",
  2516 => x"14200000",
  2517 => x"15200000",
  2518 => x"53442069",
  2519 => x"6e69742e",
  2520 => x"2e2e0a00",
  2521 => x"53442063",
  2522 => x"61726420",
  2523 => x"72657365",
  2524 => x"74206661",
  2525 => x"696c6564",
  2526 => x"210a0000",
  2527 => x"53444843",
  2528 => x"20657272",
  2529 => x"6f72210a",
  2530 => x"00000000",
  2531 => x"57726974",
  2532 => x"65206661",
  2533 => x"696c6564",
  2534 => x"0a000000",
  2535 => x"52656164",
  2536 => x"20666169",
  2537 => x"6c65640a",
  2538 => x"00000000",
  2539 => x"43617264",
  2540 => x"20696e69",
  2541 => x"74206661",
  2542 => x"696c6564",
  2543 => x"0a000000",
  2544 => x"46415431",
  2545 => x"36202020",
  2546 => x"00000000",
  2547 => x"46415433",
  2548 => x"32202020",
  2549 => x"00000000",
  2550 => x"4e6f2070",
  2551 => x"61727469",
  2552 => x"74696f6e",
  2553 => x"20736967",
  2554 => x"0a000000",
  2555 => x"42616420",
  2556 => x"70617274",
  2557 => x"0a000000",
  2558 => x"4261636b",
  2559 => x"00000000",
  2560 => x"00000002",
  2561 => x"00000000",
  2562 => x"00000010",
  2563 => x"00000002",
  2564 => x"00002584",
  2565 => x"00000a54",
  2566 => x"00000002",
  2567 => x"000025a0",
  2568 => x"00000a54",
  2569 => x"00000002",
  2570 => x"000025bc",
  2571 => x"0000037f",
  2572 => x"00000001",
  2573 => x"000025c4",
  2574 => x"00000000",
  2575 => x"00000001",
  2576 => x"000025d0",
  2577 => x"00000001",
  2578 => x"00000001",
  2579 => x"000025e0",
  2580 => x"00000002",
  2581 => x"00000002",
  2582 => x"000025f0",
  2583 => x"00002537",
  2584 => x"00000002",
  2585 => x"00002604",
  2586 => x"00002522",
  2587 => x"00000003",
  2588 => x"000028ac",
  2589 => x"00000002",
  2590 => x"00000003",
  2591 => x"0000289c",
  2592 => x"00000004",
  2593 => x"00000002",
  2594 => x"00002614",
  2595 => x"00000ffd",
  2596 => x"00000000",
  2597 => x"00000000",
  2598 => x"00000000",
  2599 => x"0000261c",
  2600 => x"00002630",
  2601 => x"00002648",
  2602 => x"00002664",
  2603 => x"00002684",
  2604 => x"0000269c",
  2605 => x"00000002",
  2606 => x"000026b4",
  2607 => x"00000a54",
  2608 => x"00000002",
  2609 => x"000025a0",
  2610 => x"00000a54",
  2611 => x"00000002",
  2612 => x"000025bc",
  2613 => x"0000037f",
  2614 => x"00000001",
  2615 => x"000025c4",
  2616 => x"00000000",
  2617 => x"00000001",
  2618 => x"000025d0",
  2619 => x"00000001",
  2620 => x"00000001",
  2621 => x"000025e0",
  2622 => x"00000002",
  2623 => x"00000002",
  2624 => x"000025f0",
  2625 => x"00002537",
  2626 => x"00000002",
  2627 => x"00002604",
  2628 => x"00002522",
  2629 => x"00000003",
  2630 => x"000028ac",
  2631 => x"00000002",
  2632 => x"00000003",
  2633 => x"0000289c",
  2634 => x"00000004",
  2635 => x"00000003",
  2636 => x"00002950",
  2637 => x"00000003",
  2638 => x"00000002",
  2639 => x"00002614",
  2640 => x"00000ffd",
  2641 => x"00000000",
  2642 => x"00000000",
  2643 => x"00000000",
  2644 => x"000026d0",
  2645 => x"000026e8",
  2646 => x"00002704",
  2647 => x"00000004",
  2648 => x"0000271c",
  2649 => x"0000295c",
  2650 => x"00000004",
  2651 => x"00002730",
  2652 => x"0000280c",
  2653 => x"00000000",
  2654 => x"00000000",
  2655 => x"00000000",
  2656 => x"00000000",
  2657 => x"00000000",
  2658 => x"00000000",
  2659 => x"00000000",
  2660 => x"00000000",
  2661 => x"00000000",
  2662 => x"00000000",
  2663 => x"00000000",
  2664 => x"00000000",
  2665 => x"00000000",
  2666 => x"00000000",
  2667 => x"00000000",
  2668 => x"00000000",
  2669 => x"00000000",
  2670 => x"00000000",
  2671 => x"00000000",
  2672 => x"00000000",
  2673 => x"00000000",
  2674 => x"00000006",
  2675 => x"00000043",
  2676 => x"00000042",
  2677 => x"0000003b",
  2678 => x"0000004b",
  2679 => x"00000033",
  2680 => x"0000001d",
  2681 => x"0000001b",
  2682 => x"0000001c",
  2683 => x"00000023",
  2684 => x"0000002b",
  2685 => x"00000000",
  2686 => x"00000000",
  2687 => x"00000002",
  2688 => x"00002e64",
  2689 => x"000022bc",
  2690 => x"00000002",
  2691 => x"00002e82",
  2692 => x"000022bc",
  2693 => x"00000002",
  2694 => x"00002ea0",
  2695 => x"000022bc",
  2696 => x"00000002",
  2697 => x"00002ebe",
  2698 => x"000022bc",
  2699 => x"00000002",
  2700 => x"00002edc",
  2701 => x"000022bc",
  2702 => x"00000002",
  2703 => x"00002efa",
  2704 => x"000022bc",
  2705 => x"00000002",
  2706 => x"00002f18",
  2707 => x"000022bc",
  2708 => x"00000002",
  2709 => x"00002f36",
  2710 => x"000022bc",
  2711 => x"00000002",
  2712 => x"00002f54",
  2713 => x"000022bc",
  2714 => x"00000002",
  2715 => x"00002f72",
  2716 => x"000022bc",
  2717 => x"00000002",
  2718 => x"00002f90",
  2719 => x"000022bc",
  2720 => x"00000002",
  2721 => x"00002fae",
  2722 => x"000022bc",
  2723 => x"00000002",
  2724 => x"00002fcc",
  2725 => x"000022bc",
  2726 => x"00000004",
  2727 => x"000027f8",
  2728 => x"00000000",
  2729 => x"00000000",
  2730 => x"00000000",
  2731 => x"00002482",
  2732 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

