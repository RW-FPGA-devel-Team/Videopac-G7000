library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sp0256_004_decoded is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sp0256_004_decoded is
	type rom is array(0 to  7775) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"18",X"12",X"00",X"2A",X"30",X"00",X"5A",X"15",X"00",X"6F",X"2F",X"00",X"9E",X"2E",X"00",
		X"CC",X"06",X"00",X"D2",X"0A",X"00",X"DC",X"16",X"00",X"F2",X"02",X"00",X"F4",X"38",X"01",X"2C",
		X"0F",X"01",X"3B",X"0A",X"01",X"45",X"08",X"01",X"4D",X"19",X"01",X"66",X"00",X"01",X"66",X"00",
		X"01",X"66",X"22",X"01",X"88",X"04",X"01",X"8C",X"00",X"01",X"8C",X"00",X"01",X"8C",X"00",X"01",
		X"8C",X"00",X"01",X"8C",X"00",X"01",X"8C",X"0D",X"01",X"99",X"25",X"01",X"BE",X"09",X"01",X"C7",
		X"03",X"01",X"CA",X"01",X"01",X"CB",X"07",X"01",X"D2",X"0F",X"01",X"E1",X"0A",X"01",X"EB",X"0D",
		X"03",X"02",X"00",X"58",X"00",X"60",X"28",X"60",X"40",X"60",X"E8",X"68",X"EC",X"12",X"90",X"75",
		X"03",X"05",X"00",X"4B",X"00",X"70",X"28",X"50",X"38",X"60",X"EC",X"68",X"F0",X"0E",X"90",X"73",
		X"03",X"05",X"00",X"40",X"00",X"60",X"28",X"50",X"40",X"70",X"F4",X"68",X"EC",X"04",X"8F",X"72",
		X"05",X"03",X"80",X"3C",X"00",X"50",X"28",X"40",X"40",X"60",X"F8",X"60",X"EC",X"04",X"97",X"61",
		X"07",X"02",X"80",X"3B",X"08",X"60",X"28",X"40",X"40",X"60",X"FC",X"60",X"EC",X"04",X"92",X"69",
		X"03",X"02",X"00",X"41",X"08",X"50",X"28",X"50",X"40",X"60",X"FC",X"68",X"EC",X"02",X"90",X"6C",
		X"05",X"02",X"80",X"4B",X"08",X"50",X"28",X"50",X"40",X"60",X"FC",X"68",X"EC",X"0A",X"93",X"67",
		X"02",X"02",X"00",X"61",X"08",X"40",X"30",X"50",X"40",X"60",X"FC",X"68",X"E8",X"0A",X"95",X"62",
		X"04",X"01",X"C0",X"6D",X"08",X"50",X"28",X"60",X"38",X"60",X"F8",X"68",X"EC",X"04",X"95",X"61",
		X"02",X"02",X"00",X"75",X"08",X"50",X"20",X"60",X"38",X"60",X"F8",X"68",X"F0",X"06",X"95",X"61",
		X"03",X"01",X"00",X"7C",X"00",X"50",X"20",X"40",X"40",X"60",X"F0",X"68",X"F0",X"02",X"95",X"63",
		X"03",X"00",X"80",X"83",X"08",X"50",X"20",X"30",X"30",X"40",X"EC",X"60",X"F4",X"F2",X"94",X"65",
		X"05",X"00",X"A0",X"7D",X"08",X"30",X"38",X"60",X"48",X"50",X"FC",X"00",X"E4",X"64",X"8E",X"6F",
		X"03",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"50",X"E8",X"02",X"0F",X"16",
		X"0A",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"10",X"34",X"5C",X"E5",X"1E",
		X"05",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"58",X"0C",X"10",X"EA",X"1F",
		X"07",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"48",X"04",X"16",X"DD",X"25",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"04",X"F8",X"00",X"D0",X"E0",X"30",X"18",X"20",X"1C",X"E8",X"18",X"04",X"00",X"00",
		X"0F",X"00",X"0C",X"72",X"30",X"D0",X"A8",X"30",X"B8",X"20",X"1C",X"E8",X"18",X"04",X"00",X"00",
		X"04",X"00",X"00",X"8B",X"30",X"D0",X"A8",X"30",X"B8",X"20",X"1C",X"E8",X"18",X"04",X"00",X"00",
		X"0F",X"03",X"80",X"1F",X"F8",X"00",X"38",X"10",X"C8",X"00",X"10",X"48",X"0C",X"D4",X"00",X"00",
		X"0B",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"80",X"2B",X"40",X"00",X"48",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"00",X"36",X"40",X"00",X"48",X"00",X"50",X"00",X"E8",X"00",X"18",X"0E",X"00",X"00",
		X"0B",X"00",X"80",X"32",X"68",X"00",X"00",X"00",X"00",X"00",X"E8",X"00",X"18",X"0E",X"00",X"00",
		X"2F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"45",X"10",X"30",X"00",X"20",X"00",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"04",X"0E",X"00",X"FF",X"20",X"30",X"98",X"20",X"20",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"03",X"00",X"00",X"FF",X"58",X"30",X"60",X"20",X"20",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"60",X"96",X"08",X"10",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"38",X"96",X"08",X"10",X"00",X"00",X"00",X"00",X"E4",X"00",X"6C",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"08",X"0C",X"3C",X"19",X"5F",X"00",X"0A",X"00",X"00",X"1E",X"C1",X"6C",X"32",
		X"03",X"00",X"28",X"46",X"F8",X"50",X"10",X"70",X"70",X"40",X"AC",X"08",X"94",X"24",X"82",X"CB",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"00",X"60",X"08",X"1C",X"00",X"40",X"00",X"00",X"08",X"18",X"60",X"AF",X"92",X"C4",X"80",
		X"0E",X"00",X"00",X"3F",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"46",X"06",X"78",X"68",X"F7",X"CF",
		X"05",X"00",X"40",X"3F",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"AC",X"06",X"E9",X"68",X"FA",X"CF",
		X"2C",X"00",X"40",X"82",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"AC",X"06",X"E9",X"68",X"FA",X"CF",
		X"0F",X"00",X"60",X"82",X"F8",X"2C",X"6C",X"66",X"38",X"1A",X"AC",X"06",X"E9",X"68",X"00",X"00",
		X"0E",X"00",X"0C",X"00",X"04",X"EA",X"8B",X"74",X"95",X"07",X"40",X"06",X"57",X"0C",X"51",X"E3",
		X"0E",X"02",X"00",X"00",X"04",X"EA",X"03",X"74",X"AD",X"07",X"40",X"06",X"57",X"0C",X"00",X"00",
		X"03",X"00",X"18",X"3E",X"6F",X"D4",X"F8",X"1F",X"CD",X"C7",X"07",X"8C",X"8C",X"00",X"02",X"11",
		X"09",X"00",X"38",X"09",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F8",X"18",X"C4",X"36",X"00",X"00",
		X"0A",X"00",X"00",X"3E",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F8",X"18",X"C4",X"36",X"00",X"00",
		X"08",X"00",X"A0",X"31",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F4",X"08",X"CC",X"42",X"00",X"00",
		X"0D",X"01",X"00",X"FC",X"D8",X"70",X"80",X"10",X"70",X"40",X"C8",X"48",X"C0",X"18",X"00",X"00",
		X"04",X"02",X"00",X"35",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"68",X"78",X"A8",X"00",X"00",
		X"09",X"03",X"80",X"2C",X"00",X"10",X"F0",X"C0",X"F0",X"D0",X"0C",X"70",X"8C",X"9E",X"00",X"00",
		X"05",X"00",X"10",X"2C",X"00",X"10",X"F0",X"C0",X"F0",X"D0",X"34",X"70",X"DC",X"9E",X"00",X"00",
		X"0D",X"00",X"14",X"90",X"F0",X"40",X"28",X"40",X"C8",X"60",X"6C",X"40",X"E0",X"5C",X"00",X"00",
		X"07",X"00",X"20",X"FD",X"F0",X"40",X"28",X"40",X"C8",X"60",X"6C",X"40",X"E0",X"5C",X"00",X"00",
		X"03",X"00",X"18",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"70",X"74",X"C0",X"00",X"00",
		X"0C",X"00",X"30",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"70",X"34",X"C0",X"00",X"00",
		X"2F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"3C",X"E2",X"9B",X"8A",X"98",X"2A",X"49",X"32",X"03",X"F0",X"8C",X"8F",X"73",X"E2",
		X"08",X"02",X"00",X"E2",X"9B",X"8A",X"98",X"2A",X"49",X"32",X"EB",X"F0",X"7C",X"8F",X"00",X"00",
		X"03",X"00",X"00",X"CD",X"0B",X"8A",X"80",X"2A",X"F1",X"32",X"EB",X"F0",X"7C",X"8F",X"00",X"00",
		X"07",X"00",X"C0",X"FA",X"10",X"10",X"00",X"60",X"C0",X"00",X"E0",X"60",X"5C",X"7E",X"00",X"00",
		X"0A",X"00",X"78",X"C4",X"A8",X"01",X"E4",X"03",X"BC",X"4F",X"03",X"C7",X"21",X"80",X"00",X"22",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"E4",X"00",X"00",X"00",
		X"07",X"00",X"00",X"3C",X"08",X"D0",X"10",X"30",X"00",X"10",X"4C",X"F8",X"00",X"F4",X"00",X"00",
		X"01",X"01",X"80",X"00",X"38",X"00",X"88",X"00",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"CE",X"38",X"00",X"88",X"00",X"E8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"A0",X"6B",X"B0",X"00",X"38",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"36",X"01",X"80",X"0E",X"D8",X"00",X"A8",X"70",X"60",X"60",X"98",X"48",X"70",X"26",X"22",X"06",
		X"08",X"01",X"00",X"0E",X"D8",X"00",X"A8",X"70",X"60",X"60",X"9C",X"48",X"78",X"26",X"3F",X"06",
		X"03",X"00",X"00",X"4E",X"D8",X"00",X"A8",X"70",X"60",X"60",X"9C",X"48",X"78",X"26",X"3F",X"06",
		X"02",X"0A",X"00",X"00",X"10",X"20",X"C8",X"00",X"F8",X"60",X"7C",X"78",X"5C",X"9A",X"02",X"9E",
		X"08",X"00",X"E8",X"C1",X"76",X"1E",X"E9",X"79",X"01",X"3F",X"04",X"00",X"DA",X"00",X"6F",X"93",
		X"0C",X"00",X"20",X"7C",X"60",X"50",X"28",X"00",X"00",X"00",X"00",X"00",X"08",X"00",X"90",X"F6",
		X"01",X"00",X"0C",X"7C",X"60",X"50",X"28",X"00",X"00",X"00",X"8C",X"00",X"84",X"00",X"1A",X"F6",
		X"03",X"0C",X"00",X"2F",X"40",X"50",X"B8",X"00",X"C0",X"00",X"8C",X"00",X"84",X"00",X"1A",X"F6",
		X"0A",X"00",X"80",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"30",X"70",X"72",X"C7",X"7C",
		X"02",X"03",X"00",X"64",X"00",X"00",X"F8",X"00",X"00",X"00",X"04",X"30",X"74",X"74",X"C7",X"7C",
		X"03",X"01",X"00",X"7C",X"00",X"50",X"20",X"40",X"40",X"60",X"F0",X"68",X"F0",X"02",X"95",X"63",
		X"03",X"00",X"80",X"83",X"08",X"50",X"20",X"30",X"30",X"40",X"EC",X"60",X"F4",X"F2",X"94",X"65",
		X"05",X"00",X"A0",X"7D",X"08",X"30",X"38",X"60",X"48",X"50",X"FC",X"00",X"E4",X"64",X"8E",X"6F",
		X"03",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"50",X"E8",X"02",X"0F",X"16",
		X"0A",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"10",X"34",X"5C",X"E5",X"1E",
		X"05",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"58",X"0C",X"10",X"EA",X"1F",
		X"07",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"48",X"04",X"16",X"DD",X"25",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"08",X"E8",X"0C",X"00",X"00",
		X"0E",X"04",X"00",X"00",X"00",X"00",X"68",X"00",X"88",X"00",X"1C",X"08",X"E8",X"0C",X"00",X"00",
		X"0F",X"03",X"80",X"1F",X"F8",X"00",X"38",X"10",X"C8",X"00",X"10",X"48",X"0C",X"D4",X"00",X"00",
		X"0B",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"80",X"2B",X"40",X"00",X"48",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"00",X"36",X"40",X"00",X"48",X"00",X"50",X"00",X"E8",X"00",X"18",X"0E",X"00",X"00",
		X"0B",X"00",X"80",X"32",X"68",X"00",X"00",X"00",X"00",X"00",X"E8",X"00",X"18",X"0E",X"00",X"00",
		X"2F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"45",X"10",X"30",X"00",X"20",X"00",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"04",X"0E",X"00",X"FF",X"20",X"30",X"98",X"20",X"20",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"03",X"00",X"00",X"FF",X"58",X"30",X"60",X"20",X"20",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"60",X"96",X"08",X"10",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"38",X"96",X"08",X"10",X"00",X"00",X"00",X"00",X"E4",X"00",X"6C",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"08",X"0C",X"3C",X"19",X"5F",X"00",X"0A",X"00",X"00",X"1E",X"C1",X"6C",X"32",
		X"03",X"00",X"28",X"46",X"F8",X"50",X"10",X"70",X"70",X"40",X"AC",X"08",X"94",X"24",X"82",X"CB",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"00",X"60",X"08",X"1C",X"00",X"40",X"00",X"00",X"08",X"18",X"60",X"AF",X"92",X"C4",X"80",
		X"0E",X"00",X"00",X"3F",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"46",X"06",X"78",X"68",X"F7",X"CF",
		X"05",X"00",X"40",X"3F",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"AC",X"06",X"E9",X"68",X"FA",X"CF",
		X"2C",X"00",X"40",X"82",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"AC",X"06",X"E9",X"68",X"FA",X"CF",
		X"0F",X"00",X"60",X"82",X"F8",X"2C",X"6C",X"66",X"38",X"1A",X"AC",X"06",X"E9",X"68",X"00",X"00",
		X"0E",X"00",X"0C",X"00",X"04",X"EA",X"8B",X"74",X"95",X"07",X"40",X"06",X"57",X"0C",X"51",X"E3",
		X"0E",X"02",X"00",X"00",X"04",X"EA",X"03",X"74",X"AD",X"07",X"40",X"06",X"57",X"0C",X"00",X"00",
		X"03",X"00",X"18",X"3E",X"6F",X"D4",X"F8",X"1F",X"CD",X"C7",X"07",X"8C",X"8C",X"00",X"02",X"11",
		X"09",X"00",X"38",X"09",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F8",X"18",X"C4",X"36",X"00",X"00",
		X"0A",X"00",X"00",X"3E",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F8",X"18",X"C4",X"36",X"00",X"00",
		X"08",X"00",X"A0",X"31",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F4",X"08",X"CC",X"42",X"00",X"00",
		X"0D",X"01",X"00",X"FC",X"D8",X"70",X"80",X"10",X"70",X"40",X"C8",X"48",X"C0",X"18",X"00",X"00",
		X"04",X"02",X"00",X"35",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"68",X"78",X"A8",X"00",X"00",
		X"09",X"03",X"80",X"2C",X"00",X"10",X"F0",X"C0",X"F0",X"D0",X"0C",X"70",X"8C",X"9E",X"00",X"00",
		X"05",X"00",X"10",X"2C",X"00",X"10",X"F0",X"C0",X"F0",X"D0",X"34",X"70",X"DC",X"9E",X"00",X"00",
		X"0D",X"00",X"14",X"90",X"F0",X"40",X"28",X"40",X"C8",X"60",X"6C",X"40",X"E0",X"5C",X"00",X"00",
		X"07",X"00",X"20",X"FD",X"F0",X"40",X"28",X"40",X"C8",X"60",X"6C",X"40",X"E0",X"5C",X"00",X"00",
		X"03",X"00",X"18",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"70",X"74",X"C0",X"00",X"00",
		X"0C",X"00",X"30",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"70",X"34",X"C0",X"00",X"00",
		X"2F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"3C",X"E2",X"9B",X"8A",X"98",X"2A",X"49",X"32",X"03",X"F0",X"8C",X"8F",X"73",X"E2",
		X"08",X"02",X"00",X"E2",X"9B",X"8A",X"98",X"2A",X"49",X"32",X"EB",X"F0",X"7C",X"8F",X"00",X"00",
		X"03",X"00",X"00",X"CD",X"0B",X"8A",X"80",X"2A",X"F1",X"32",X"EB",X"F0",X"7C",X"8F",X"00",X"00",
		X"07",X"00",X"C0",X"FA",X"10",X"10",X"00",X"60",X"C0",X"00",X"E0",X"60",X"5C",X"7E",X"00",X"00",
		X"0A",X"00",X"78",X"C4",X"A8",X"01",X"E4",X"03",X"BC",X"4F",X"03",X"C7",X"21",X"80",X"00",X"22",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"E4",X"00",X"00",X"00",
		X"07",X"00",X"00",X"3C",X"08",X"D0",X"10",X"30",X"00",X"10",X"4C",X"F8",X"00",X"F4",X"00",X"00",
		X"06",X"00",X"C0",X"E9",X"00",X"00",X"68",X"00",X"88",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"03",X"80",X"1F",X"F8",X"00",X"38",X"10",X"C8",X"00",X"10",X"48",X"0C",X"D4",X"00",X"00",
		X"0B",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"80",X"2B",X"40",X"00",X"48",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"00",X"36",X"40",X"00",X"48",X"00",X"50",X"00",X"E8",X"00",X"18",X"0E",X"00",X"00",
		X"0B",X"00",X"80",X"32",X"68",X"00",X"00",X"00",X"00",X"00",X"E8",X"00",X"18",X"0E",X"00",X"00",
		X"2F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"45",X"10",X"30",X"00",X"20",X"00",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"04",X"0E",X"00",X"FF",X"20",X"30",X"98",X"20",X"20",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"03",X"00",X"00",X"FF",X"58",X"30",X"60",X"20",X"20",X"00",X"08",X"00",X"0C",X"F0",X"00",X"00",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"97",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"60",X"96",X"08",X"10",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"38",X"96",X"08",X"10",X"00",X"00",X"00",X"00",X"E4",X"00",X"6C",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"08",X"0C",X"3C",X"19",X"5F",X"00",X"0A",X"00",X"00",X"1E",X"C1",X"6C",X"32",
		X"03",X"00",X"28",X"46",X"F8",X"50",X"10",X"70",X"70",X"40",X"AC",X"08",X"94",X"24",X"82",X"CB",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"38",X"00",X"60",X"08",X"1C",X"00",X"40",X"00",X"00",X"08",X"18",X"60",X"AF",X"92",X"C4",X"80",
		X"0E",X"00",X"00",X"3F",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"46",X"06",X"78",X"68",X"F7",X"CF",
		X"05",X"00",X"40",X"3F",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"AC",X"06",X"E9",X"68",X"FA",X"CF",
		X"2C",X"00",X"40",X"82",X"94",X"2C",X"C0",X"66",X"60",X"1A",X"AC",X"06",X"E9",X"68",X"FA",X"CF",
		X"0F",X"00",X"60",X"82",X"F8",X"2C",X"6C",X"66",X"38",X"1A",X"AC",X"06",X"E9",X"68",X"00",X"00",
		X"0E",X"00",X"0C",X"00",X"04",X"EA",X"8B",X"74",X"95",X"07",X"40",X"06",X"57",X"0C",X"51",X"E3",
		X"0E",X"02",X"00",X"00",X"04",X"EA",X"03",X"74",X"AD",X"07",X"40",X"06",X"57",X"0C",X"00",X"00",
		X"03",X"00",X"18",X"3E",X"6F",X"D4",X"F8",X"1F",X"CD",X"C7",X"07",X"8C",X"8C",X"00",X"02",X"11",
		X"09",X"00",X"38",X"09",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F8",X"18",X"C4",X"36",X"00",X"00",
		X"0A",X"00",X"00",X"3E",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F8",X"18",X"C4",X"36",X"00",X"00",
		X"08",X"00",X"A0",X"31",X"B0",X"70",X"08",X"50",X"A8",X"50",X"F4",X"08",X"CC",X"42",X"00",X"00",
		X"0D",X"01",X"00",X"FC",X"D8",X"70",X"80",X"10",X"70",X"40",X"C8",X"48",X"C0",X"18",X"00",X"00",
		X"04",X"02",X"00",X"35",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"68",X"78",X"A8",X"00",X"00",
		X"09",X"03",X"80",X"2C",X"00",X"10",X"F0",X"C0",X"F0",X"D0",X"0C",X"70",X"8C",X"9E",X"00",X"00",
		X"05",X"00",X"10",X"2C",X"00",X"10",X"F0",X"C0",X"F0",X"D0",X"34",X"70",X"DC",X"9E",X"00",X"00",
		X"0D",X"00",X"14",X"90",X"F0",X"40",X"28",X"40",X"C8",X"60",X"6C",X"40",X"E0",X"5C",X"00",X"00",
		X"07",X"00",X"20",X"FD",X"F0",X"40",X"28",X"40",X"C8",X"60",X"6C",X"40",X"E0",X"5C",X"00",X"00",
		X"03",X"00",X"18",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"9C",X"70",X"74",X"C0",X"00",X"00",
		X"0C",X"00",X"30",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"4C",X"70",X"34",X"C0",X"00",X"00",
		X"2F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"3C",X"E2",X"9B",X"8A",X"98",X"2A",X"49",X"32",X"03",X"F0",X"8C",X"8F",X"73",X"E2",
		X"08",X"02",X"00",X"E2",X"9B",X"8A",X"98",X"2A",X"49",X"32",X"EB",X"F0",X"7C",X"8F",X"00",X"00",
		X"03",X"00",X"00",X"CD",X"0B",X"8A",X"80",X"2A",X"F1",X"32",X"EB",X"F0",X"7C",X"8F",X"00",X"00",
		X"07",X"00",X"C0",X"FA",X"10",X"10",X"00",X"60",X"C0",X"00",X"E0",X"60",X"5C",X"7E",X"00",X"00",
		X"0A",X"00",X"78",X"C4",X"A8",X"01",X"E4",X"03",X"BC",X"4F",X"03",X"C7",X"21",X"80",X"00",X"22",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"80",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"00",X"E4",X"00",X"00",X"00",
		X"07",X"00",X"00",X"3C",X"08",X"D0",X"10",X"30",X"00",X"10",X"4C",X"F8",X"00",X"F4",X"00",X"00",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"40",X"40",X"98",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"1A",X"92",X"F3",X"A6",X"37",X"E2",X"69",X"21",X"50",X"15",X"49",X"C8",X"98",X"DA",
		X"0E",X"0C",X"00",X"9B",X"F8",X"00",X"B0",X"00",X"08",X"30",X"78",X"00",X"90",X"60",X"00",X"00",
		X"08",X"00",X"F0",X"0B",X"90",X"20",X"C2",X"3F",X"83",X"ED",X"80",X"84",X"26",X"08",X"40",X"0D",
		X"0E",X"00",X"A0",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"A8",X"60",X"24",X"FC",X"00",X"00",
		X"16",X"00",X"20",X"86",X"18",X"20",X"A0",X"30",X"F8",X"60",X"80",X"58",X"B0",X"5C",X"CA",X"4A",
		X"05",X"00",X"04",X"86",X"18",X"20",X"A0",X"30",X"F8",X"60",X"E4",X"58",X"E0",X"5C",X"F8",X"4A",
		X"0E",X"00",X"0F",X"24",X"01",X"0B",X"00",X"38",X"00",X"88",X"86",X"60",X"2B",X"E4",X"31",X"20",
		X"0F",X"00",X"54",X"CE",X"83",X"70",X"23",X"0D",X"BC",X"34",X"FB",X"E7",X"CA",X"32",X"AE",X"9A",
		X"07",X"00",X"08",X"F8",X"2B",X"70",X"5B",X"0D",X"F4",X"34",X"FB",X"E7",X"CA",X"32",X"AE",X"9A",
		X"07",X"00",X"1C",X"47",X"00",X"60",X"00",X"00",X"70",X"50",X"80",X"10",X"88",X"DC",X"95",X"07",
		X"07",X"00",X"C0",X"47",X"38",X"60",X"50",X"00",X"F0",X"50",X"80",X"10",X"88",X"DC",X"95",X"07",
		X"02",X"01",X"80",X"47",X"28",X"60",X"48",X"20",X"D0",X"50",X"8C",X"10",X"A4",X"D4",X"92",X"0F",
		X"07",X"01",X"40",X"47",X"28",X"60",X"48",X"20",X"D0",X"50",X"88",X"00",X"9C",X"DA",X"85",X"15",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"26",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"01",X"00",X"40",X"A8",X"00",X"20",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"20",X"22",X"A8",X"00",X"20",X"00",X"08",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"14",X"88",X"D0",X"38",X"C0",X"10",X"F0",X"1C",X"00",X"00",X"00",X"FC",X"00",
		X"0C",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"01",X"80",X"FC",X"08",X"00",X"10",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"78",X"63",X"50",X"FF",X"F8",X"90",X"7F",X"F0",X"EB",X"E0",X"67",X"1A",X"28",X"76",
		X"03",X"02",X"80",X"4F",X"A0",X"FF",X"F8",X"90",X"E7",X"F0",X"EB",X"E0",X"67",X"1A",X"28",X"76",
		X"04",X"01",X"C0",X"B1",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"28",X"98",X"FE",X"6D",X"18",
		X"0E",X"00",X"00",X"5F",X"D0",X"30",X"98",X"40",X"A8",X"10",X"3C",X"48",X"98",X"00",X"E8",X"F4",
		X"0E",X"05",X"00",X"5F",X"D0",X"30",X"98",X"40",X"A8",X"10",X"F0",X"48",X"70",X"00",X"52",X"F4",
		X"09",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"14",X"0E",X"00",X"83",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"60",X"80",X"FA",X"00",X"00",
		X"03",X"00",X"00",X"CC",X"B0",X"40",X"78",X"60",X"E8",X"60",X"84",X"70",X"F4",X"90",X"00",X"00",
		X"04",X"06",X"C0",X"A7",X"39",X"4C",X"EE",X"D8",X"C4",X"41",X"C0",X"36",X"0B",X"3F",X"07",X"8D",
		X"08",X"01",X"00",X"DA",X"D1",X"4C",X"E6",X"D8",X"DC",X"41",X"C0",X"36",X"0B",X"3F",X"00",X"00",
		X"01",X"00",X"20",X"AF",X"80",X"00",X"C0",X"30",X"C8",X"40",X"A4",X"18",X"48",X"C2",X"00",X"00",
		X"07",X"00",X"00",X"D3",X"80",X"00",X"C0",X"30",X"C8",X"40",X"A4",X"18",X"48",X"C2",X"00",X"00",
		X"0D",X"00",X"20",X"94",X"80",X"00",X"C0",X"30",X"C8",X"40",X"A4",X"18",X"48",X"C2",X"00",X"00",
		X"05",X"00",X"A0",X"7D",X"08",X"30",X"38",X"60",X"48",X"50",X"FC",X"00",X"E4",X"64",X"00",X"00",
		X"0F",X"00",X"30",X"7D",X"08",X"30",X"38",X"60",X"48",X"50",X"38",X"00",X"C8",X"64",X"00",X"00",
		X"0F",X"03",X"00",X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",
		X"08",X"00",X"1C",X"00",X"20",X"00",X"30",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"0A",X"00",X"DB",X"00",X"70",X"F8",X"60",X"70",X"10",X"CC",X"18",X"00",X"F0",X"00",X"00",
		X"01",X"00",X"08",X"01",X"60",X"00",X"88",X"00",X"A0",X"40",X"48",X"38",X"6C",X"70",X"00",X"00",
		X"03",X"01",X"80",X"E3",X"68",X"70",X"E0",X"20",X"B0",X"30",X"3C",X"20",X"3C",X"A0",X"00",X"00",
		X"04",X"01",X"C0",X"D9",X"68",X"80",X"E8",X"40",X"98",X"40",X"1C",X"18",X"38",X"90",X"00",X"00",
		X"02",X"00",X"E0",X"E8",X"58",X"B0",X"E0",X"40",X"88",X"70",X"08",X"18",X"24",X"9E",X"00",X"00",
		X"0C",X"00",X"00",X"C1",X"18",X"60",X"80",X"50",X"D8",X"30",X"94",X"08",X"D8",X"66",X"00",X"00",
		X"07",X"00",X"20",X"C0",X"F8",X"40",X"70",X"10",X"D8",X"60",X"84",X"00",X"D8",X"70",X"00",X"00",
		X"0E",X"00",X"20",X"A0",X"F8",X"40",X"70",X"10",X"D8",X"60",X"84",X"00",X"D8",X"70",X"00",X"00",
		X"04",X"06",X"00",X"46",X"F8",X"50",X"20",X"60",X"38",X"60",X"E4",X"60",X"EC",X"FE",X"00",X"00",
		X"01",X"01",X"00",X"46",X"B0",X"50",X"30",X"60",X"70",X"60",X"E4",X"60",X"EC",X"FE",X"00",X"00",
		X"03",X"04",X"00",X"3D",X"16",X"8A",X"F0",X"17",X"A8",X"55",X"DF",X"37",X"F9",X"4F",X"11",X"04",
		X"0F",X"0C",X"00",X"45",X"16",X"8A",X"F0",X"17",X"A8",X"55",X"CF",X"17",X"E9",X"4B",X"11",X"04",
		X"0E",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"18",X"51",X"08",X"50",X"78",X"30",X"90",X"10",X"00",X"10",X"28",X"80",X"00",X"00",
		X"0F",X"02",X"00",X"51",X"E8",X"50",X"88",X"30",X"38",X"10",X"00",X"10",X"28",X"80",X"00",X"00",
		X"04",X"01",X"C0",X"51",X"B0",X"50",X"30",X"30",X"E8",X"10",X"00",X"10",X"28",X"80",X"00",X"00",
		X"06",X"00",X"40",X"4D",X"C0",X"80",X"38",X"F0",X"E8",X"D0",X"E4",X"28",X"24",X"7E",X"00",X"00",
		X"01",X"00",X"70",X"9F",X"98",X"80",X"88",X"F0",X"B8",X"D0",X"E4",X"28",X"24",X"7E",X"00",X"00",
		X"0C",X"00",X"20",X"99",X"98",X"B0",X"90",X"20",X"B0",X"00",X"F4",X"20",X"04",X"86",X"00",X"00",
		X"05",X"00",X"20",X"73",X"98",X"B0",X"90",X"20",X"B0",X"00",X"F4",X"20",X"04",X"86",X"00",X"00",
		X"06",X"00",X"28",X"78",X"98",X"B0",X"90",X"20",X"B0",X"00",X"F0",X"00",X"10",X"86",X"00",X"00",
		X"27",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"80",X"EC",X"18",X"00",X"90",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"80",X"E8",X"18",X"00",X"90",X"00",X"F0",X"00",X"04",X"E0",X"FC",X"0E",X"00",X"00",
		X"0F",X"00",X"00",X"8F",X"F0",X"00",X"60",X"00",X"C8",X"00",X"04",X"E0",X"FC",X"0E",X"00",X"00",
		X"0C",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"04",X"00",X"3C",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"E0",X"08",X"FE",X"00",X"00",
		X"0A",X"00",X"00",X"2D",X"E0",X"E0",X"00",X"10",X"E8",X"E0",X"E8",X"C0",X"20",X"00",X"00",X"00",
		X"04",X"00",X"20",X"20",X"A8",X"70",X"A8",X"10",X"A0",X"10",X"D0",X"30",X"58",X"32",X"00",X"00",
		X"0E",X"02",X"00",X"33",X"D8",X"00",X"98",X"40",X"38",X"50",X"0C",X"00",X"64",X"5C",X"00",X"00",
		X"0E",X"00",X"60",X"09",X"28",X"20",X"20",X"20",X"F0",X"60",X"94",X"78",X"4C",X"34",X"00",X"00",
		X"06",X"08",X"00",X"23",X"78",X"20",X"00",X"20",X"00",X"60",X"94",X"78",X"4C",X"34",X"00",X"00",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"03",X"00",X"40",X"40",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"02",X"00",X"33",X"50",X"F0",X"78",X"10",X"F0",X"E0",X"F0",X"18",X"00",X"06",X"00",X"00",
		X"06",X"04",X"00",X"8C",X"68",X"10",X"E8",X"00",X"E0",X"00",X"AC",X"10",X"60",X"E0",X"00",X"00",
		X"0E",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"36",X"00",X"10",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"66",X"81",X"C0",X"59",X"0F",
		X"0A",X"01",X"80",X"AF",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"66",X"81",X"C0",X"59",X"0F",
		X"01",X"01",X"40",X"A2",X"20",X"00",X"60",X"00",X"14",X"00",X"02",X"66",X"81",X"C0",X"59",X"0F",
		X"09",X"00",X"18",X"A2",X"20",X"00",X"60",X"00",X"14",X"00",X"1E",X"66",X"00",X"C0",X"C0",X"0F",
		X"09",X"0C",X"00",X"AF",X"20",X"00",X"60",X"00",X"14",X"00",X"3C",X"5E",X"F0",X"CE",X"B5",X"15",
		X"0C",X"00",X"00",X"C1",X"8C",X"6C",X"70",X"66",X"D8",X"7A",X"44",X"0C",X"F0",X"66",X"E1",X"1F",
		X"06",X"00",X"10",X"C1",X"8C",X"6C",X"70",X"66",X"D8",X"7A",X"9C",X"0C",X"29",X"66",X"D9",X"1F",
		X"0A",X"04",X"00",X"11",X"24",X"3E",X"DC",X"62",X"F8",X"18",X"EC",X"18",X"00",X"AD",X"16",X"0F",
		X"0E",X"00",X"1C",X"11",X"24",X"3E",X"DC",X"62",X"F8",X"18",X"CA",X"18",X"99",X"AD",X"00",X"00",
		X"0D",X"00",X"80",X"7E",X"24",X"3E",X"DC",X"62",X"F8",X"18",X"CA",X"18",X"99",X"AD",X"00",X"00",
		X"03",X"01",X"C0",X"7F",X"1C",X"4C",X"DC",X"66",X"E4",X"16",X"CA",X"10",X"93",X"B7",X"00",X"00",
		X"0E",X"00",X"30",X"7C",X"1C",X"4C",X"DC",X"66",X"E4",X"16",X"CA",X"10",X"93",X"B7",X"00",X"00",
		X"08",X"0E",X"00",X"BF",X"94",X"0E",X"D4",X"54",X"18",X"70",X"7A",X"08",X"A2",X"8F",X"00",X"00",
		X"05",X"00",X"14",X"F0",X"54",X"0E",X"84",X"54",X"E8",X"70",X"7A",X"08",X"A2",X"8F",X"00",X"00",
		X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"0E",X"00",X"44",X"E0",X"F0",X"FC",X"00",X"00",X"FC",X"1E",X"00",X"FD",X"0A",X"00",X"00",
		X"04",X"00",X"14",X"3E",X"E0",X"F0",X"FC",X"00",X"00",X"FC",X"02",X"FA",X"FB",X"14",X"00",X"00",
		X"09",X"00",X"02",X"96",X"C1",X"FF",X"E7",X"D7",X"97",X"8C",X"4E",X"56",X"C3",X"D1",X"9F",X"B2",
		X"04",X"06",X"C0",X"86",X"F1",X"D6",X"F1",X"37",X"7A",X"59",X"4F",X"A0",X"DA",X"B5",X"3D",X"B8",
		X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"0A",X"00",X"A8",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"60",X"00",X"EE",X"00",X"00",
		X"04",X"00",X"60",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"60",X"00",X"EE",X"00",X"00",
		X"0B",X"00",X"80",X"86",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"60",X"88",X"EE",X"00",X"00",
		X"0F",X"00",X"C0",X"9E",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"60",X"88",X"EE",X"00",X"00",
		X"0C",X"00",X"80",X"9E",X"00",X"00",X"00",X"00",X"00",X"00",X"08",X"40",X"68",X"EC",X"00",X"00",
		X"0F",X"00",X"28",X"A4",X"78",X"00",X"C0",X"00",X"80",X"00",X"08",X"40",X"68",X"EC",X"00",X"00",
		X"03",X"04",X"00",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"B4",X"48",X"1C",X"B2",X"00",X"00",
		X"09",X"02",X"00",X"4F",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"48",X"88",X"B2",X"00",X"00",
		X"03",X"00",X"00",X"C3",X"E8",X"00",X"B8",X"00",X"F8",X"00",X"20",X"48",X"88",X"B2",X"00",X"00",
		X"03",X"00",X"1C",X"69",X"18",X"40",X"A0",X"60",X"80",X"10",X"80",X"68",X"A4",X"8C",X"00",X"00",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"0C",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"FC",X"E8",X"E4",X"02",X"00",X"00",
		X"13",X"0E",X"00",X"0D",X"E0",X"00",X"48",X"00",X"90",X"00",X"FC",X"E8",X"E4",X"02",X"00",X"00",
		X"02",X"05",X"00",X"39",X"F6",X"64",X"E8",X"0D",X"BE",X"3A",X"AD",X"35",X"7D",X"54",X"0F",X"87",
		X"03",X"0E",X"00",X"7F",X"3E",X"64",X"28",X"0D",X"B6",X"3A",X"AD",X"35",X"7D",X"54",X"00",X"00",
		X"0B",X"01",X"C0",X"7F",X"FE",X"64",X"58",X"0D",X"96",X"3A",X"AD",X"35",X"7D",X"54",X"00",X"00",
		X"0E",X"02",X"00",X"78",X"E6",X"94",X"70",X"2D",X"9E",X"4A",X"AD",X"35",X"8D",X"52",X"00",X"00",
		X"03",X"06",X"00",X"E9",X"E6",X"94",X"70",X"2D",X"9E",X"4A",X"AD",X"35",X"8D",X"52",X"00",X"00",
		X"0F",X"00",X"08",X"E9",X"7E",X"94",X"B0",X"2D",X"AE",X"4A",X"AD",X"35",X"8D",X"52",X"00",X"00",
		X"09",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"04",X"00",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"E8",X"E0",X"0C",X"00",X"00",
		X"0E",X"00",X"00",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"E8",X"E0",X"0C",X"00",X"00",
		X"02",X"00",X"60",X"7E",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"20",X"B6",X"00",X"00",
		X"01",X"08",X"00",X"00",X"F0",X"00",X"58",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"01",X"00",X"00",X"F0",X"00",X"58",X"00",X"40",X"00",X"1C",X"00",X"9C",X"00",X"00",X"00",
		X"0E",X"02",X"00",X"D7",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"08",X"8C",X"28",X"00",X"00",
		X"09",X"00",X"00",X"CE",X"0C",X"08",X"F8",X"FE",X"18",X"02",X"70",X"0A",X"89",X"2C",X"0A",X"F1",
		X"0D",X"01",X"80",X"CD",X"10",X"0C",X"DC",X"FA",X"00",X"FC",X"6E",X"FC",X"93",X"2A",X"0A",X"F1",
		X"03",X"00",X"28",X"43",X"10",X"0C",X"DC",X"FA",X"00",X"FC",X"6E",X"FC",X"93",X"2A",X"0A",X"F1",
		X"0F",X"01",X"00",X"0A",X"14",X"40",X"C8",X"62",X"24",X"1E",X"16",X"30",X"00",X"A1",X"00",X"00",
		X"08",X"00",X"10",X"31",X"04",X"38",X"C4",X"74",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1B",X"00",X"38",X"09",X"B0",X"00",X"28",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"43",X"B0",X"00",X"28",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0C",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"20",X"96",X"80",X"60",X"B0",X"60",X"10",X"20",X"38",X"00",X"20",X"D4",X"00",X"00",
		X"02",X"02",X"00",X"E1",X"28",X"60",X"68",X"60",X"60",X"20",X"38",X"00",X"20",X"D4",X"00",X"00",
		X"08",X"00",X"00",X"60",X"28",X"60",X"68",X"60",X"60",X"20",X"38",X"00",X"20",X"D4",X"00",X"00",
		X"05",X"00",X"40",X"4D",X"D8",X"60",X"28",X"60",X"A8",X"20",X"38",X"00",X"20",X"D4",X"00",X"00",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"08",X"00",X"40",X"B3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"18",X"5C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"20",X"4A",X"B8",X"00",X"38",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"30",X"4D",X"B8",X"00",X"38",X"00",X"80",X"00",X"E8",X"F8",X"E0",X"FE",X"00",X"00",
		X"03",X"00",X"10",X"35",X"B8",X"40",X"20",X"70",X"E8",X"40",X"88",X"28",X"34",X"AC",X"00",X"00",
		X"03",X"00",X"10",X"26",X"B8",X"40",X"20",X"70",X"E8",X"40",X"A0",X"28",X"14",X"B4",X"00",X"00",
		X"0A",X"00",X"00",X"1C",X"40",X"70",X"70",X"70",X"A0",X"60",X"8C",X"60",X"EC",X"F4",X"00",X"00",
		X"03",X"00",X"40",X"1C",X"30",X"70",X"78",X"70",X"00",X"60",X"8C",X"60",X"EC",X"F4",X"00",X"00",
		X"0A",X"00",X"70",X"29",X"30",X"70",X"78",X"70",X"00",X"60",X"A4",X"40",X"EC",X"EE",X"00",X"00",
		X"0D",X"01",X"80",X"29",X"18",X"70",X"E0",X"70",X"90",X"60",X"A4",X"40",X"EC",X"EE",X"00",X"00",
		X"0E",X"03",X"80",X"29",X"20",X"70",X"94",X"70",X"98",X"60",X"A4",X"40",X"EC",X"EE",X"00",X"00",
		X"06",X"00",X"10",X"0F",X"B0",X"08",X"E4",X"12",X"E4",X"3A",X"8A",X"1C",X"E6",X"D5",X"4A",X"75",
		X"0C",X"00",X"10",X"0F",X"B0",X"08",X"E4",X"12",X"E4",X"3A",X"88",X"28",X"E6",X"DD",X"3B",X"75",
		X"03",X"00",X"04",X"0F",X"80",X"08",X"E0",X"12",X"B4",X"3A",X"88",X"28",X"E6",X"DD",X"3B",X"75",
		X"08",X"00",X"C0",X"09",X"80",X"08",X"E8",X"12",X"94",X"3A",X"88",X"28",X"E6",X"DD",X"3B",X"75",
		X"08",X"00",X"C0",X"FD",X"80",X"0A",X"D8",X"0A",X"78",X"30",X"88",X"28",X"ED",X"EB",X"3C",X"78",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"84",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"0C",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"38",X"90",X"00",X"00",X"50",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"CA",X"00",X"00",X"50",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"80",X"7D",X"08",X"50",X"28",X"50",X"18",X"10",X"BC",X"58",X"08",X"FA",X"00",X"00",
		X"08",X"00",X"C0",X"7D",X"50",X"50",X"30",X"50",X"B0",X"10",X"BC",X"58",X"08",X"FA",X"00",X"00",
		X"18",X"06",X"00",X"09",X"20",X"00",X"00",X"40",X"80",X"30",X"9C",X"48",X"A8",X"32",X"21",X"1F",
		X"04",X"02",X"00",X"F0",X"30",X"20",X"C0",X"60",X"F0",X"10",X"00",X"00",X"CC",X"18",X"57",X"D8",
		X"09",X"00",X"28",X"E2",X"B0",X"30",X"70",X"20",X"B8",X"40",X"B0",X"58",X"F8",X"CC",X"01",X"56",
		X"03",X"00",X"1C",X"F1",X"B0",X"30",X"70",X"20",X"B8",X"40",X"B8",X"60",X"04",X"CA",X"09",X"49",
		X"09",X"00",X"04",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"60",X"C0",X"04",X"3F",X"06",
		X"02",X"0A",X"00",X"1C",X"00",X"00",X"08",X"10",X"00",X"00",X"3C",X"60",X"C0",X"02",X"42",X"08",
		X"04",X"07",X"00",X"7F",X"00",X"50",X"20",X"30",X"40",X"60",X"E8",X"58",X"EC",X"0C",X"AD",X"67",
		X"01",X"01",X"C0",X"A1",X"08",X"50",X"10",X"20",X"40",X"70",X"E4",X"60",X"AC",X"5C",X"E7",X"0B",
		X"08",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"18",X"48",X"F4",X"F6",X"EB",X"2E",
		X"07",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"58",X"00",X"08",X"EC",X"20",
		X"0D",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"50",X"10",X"1C",X"EB",X"30",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"3C",X"50",X"10",X"24",X"E5",X"2B",
		X"06",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"48",X"0C",X"2E",X"D6",X"21",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"07",X"00",X"28",X"08",X"50",X"20",X"40",X"38",X"50",X"F0",X"60",X"E0",X"14",X"AB",X"57",
		X"05",X"06",X"00",X"3C",X"08",X"50",X"18",X"30",X"38",X"50",X"F0",X"58",X"B0",X"52",X"DD",X"15",
		X"06",X"05",X"00",X"3D",X"08",X"50",X"18",X"20",X"38",X"40",X"F0",X"58",X"E0",X"14",X"AF",X"51",
		X"05",X"05",X"00",X"3A",X"08",X"50",X"18",X"30",X"38",X"50",X"F0",X"60",X"E0",X"16",X"AC",X"56",
		X"05",X"03",X"00",X"39",X"08",X"40",X"10",X"30",X"38",X"50",X"EC",X"60",X"E0",X"0A",X"AD",X"59",
		X"04",X"00",X"C0",X"3B",X"00",X"00",X"10",X"30",X"40",X"60",X"F0",X"28",X"E4",X"42",X"99",X"5C",
		X"05",X"01",X"C0",X"42",X"00",X"50",X"38",X"50",X"40",X"60",X"E8",X"40",X"E8",X"14",X"A2",X"50",
		X"02",X"04",X"00",X"52",X"08",X"60",X"20",X"40",X"40",X"70",X"EC",X"60",X"E4",X"0E",X"AD",X"47",
		X"04",X"01",X"80",X"6E",X"08",X"60",X"20",X"40",X"38",X"50",X"F0",X"68",X"DC",X"10",X"AE",X"46",
		X"03",X"01",X"40",X"94",X"08",X"50",X"20",X"40",X"38",X"60",X"F4",X"58",X"E8",X"04",X"A0",X"5B",
		X"03",X"01",X"C0",X"95",X"08",X"50",X"20",X"50",X"30",X"40",X"F8",X"60",X"F4",X"0C",X"92",X"72",
		X"02",X"01",X"80",X"9D",X"08",X"50",X"20",X"50",X"38",X"60",X"F8",X"58",X"F0",X"0E",X"99",X"62",
		X"02",X"00",X"E0",X"9C",X"08",X"50",X"28",X"50",X"40",X"60",X"FC",X"60",X"E8",X"0A",X"9E",X"5B",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"AC",X"18",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"04",X"38",X"18",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"38",X"18",X"00",X"20",X"00",X"00",X"00",X"80",X"00",X"CC",X"00",X"00",X"00",
		X"0E",X"0E",X"00",X"07",X"C0",X"00",X"D8",X"00",X"E8",X"00",X"80",X"00",X"CC",X"00",X"00",X"00",
		X"0A",X"00",X"18",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"F4",X"F8",X"0C",X"02",X"00",X"00",
		X"08",X"02",X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"18",X"9C",X"42",X"00",X"00",
		X"03",X"0E",X"00",X"75",X"F8",X"30",X"E0",X"30",X"00",X"10",X"30",X"00",X"B8",X"3A",X"00",X"00",
		X"06",X"03",X"80",X"75",X"80",X"30",X"E0",X"30",X"08",X"10",X"30",X"00",X"B8",X"3A",X"00",X"00",
		X"35",X"00",X"20",X"F7",X"48",X"30",X"08",X"30",X"40",X"10",X"30",X"00",X"B8",X"3A",X"00",X"00",
		X"02",X"04",X"00",X"F7",X"48",X"30",X"08",X"30",X"40",X"10",X"C8",X"00",X"7C",X"3A",X"C0",X"00",
		X"03",X"00",X"80",X"AD",X"E0",X"30",X"50",X"30",X"00",X"10",X"C8",X"00",X"7C",X"3A",X"C0",X"00",
		X"04",X"0E",X"00",X"9D",X"60",X"30",X"30",X"30",X"78",X"10",X"C8",X"00",X"7C",X"3A",X"C0",X"00",
		X"02",X"01",X"10",X"23",X"29",X"EB",X"09",X"F2",X"4D",X"31",X"44",X"BB",X"61",X"A0",X"BC",X"44",
		X"0A",X"01",X"40",X"C6",X"C0",X"40",X"E0",X"20",X"60",X"70",X"7C",X"40",X"34",X"DC",X"98",X"5F",
		X"0D",X"01",X"80",X"B9",X"D8",X"10",X"C8",X"30",X"70",X"70",X"5C",X"50",X"18",X"DA",X"A7",X"52",
		X"0E",X"00",X"50",X"E7",X"20",X"10",X"E8",X"30",X"68",X"70",X"5C",X"50",X"18",X"DA",X"A7",X"52",
		X"0F",X"00",X"08",X"80",X"20",X"10",X"E8",X"30",X"68",X"70",X"5C",X"50",X"18",X"DA",X"A7",X"52",
		X"0D",X"0C",X"00",X"AC",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"70",X"84",X"E4",X"00",X"00",
		X"0D",X"04",X"80",X"EC",X"05",X"3E",X"46",X"24",X"1F",X"CB",X"28",X"F0",X"CA",X"D7",X"00",X"15",
		X"20",X"0C",X"00",X"EF",X"00",X"00",X"00",X"00",X"00",X"00",X"98",X"20",X"58",X"F2",X"00",X"00",
		X"04",X"00",X"00",X"EF",X"40",X"00",X"70",X"00",X"20",X"00",X"98",X"20",X"58",X"F2",X"00",X"00",
		X"07",X"00",X"00",X"A4",X"F3",X"08",X"DE",X"C1",X"4A",X"45",X"DF",X"53",X"73",X"F4",X"F1",X"14",
		X"0D",X"01",X"C0",X"DF",X"13",X"08",X"5E",X"C1",X"7A",X"45",X"DF",X"53",X"73",X"F4",X"00",X"00",
		X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"04",X"00",X"ED",X"9C",X"2E",X"74",X"50",X"E4",X"5A",X"4C",X"08",X"07",X"3F",X"DA",X"D1",
		X"09",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"02",X"C0",X"F2",X"90",X"1E",X"81",X"04",X"1F",X"7B",X"5C",X"64",X"7E",X"BA",X"9E",X"92",
		X"0C",X"00",X"50",X"B2",X"50",X"66",X"60",X"44",X"B0",X"7E",X"64",X"50",X"FE",X"EF",X"24",X"BE",
		X"0B",X"02",X"00",X"B2",X"04",X"66",X"00",X"44",X"70",X"7E",X"64",X"50",X"FE",X"EF",X"24",X"BE",
		X"03",X"00",X"80",X"15",X"51",X"CC",X"00",X"0A",X"0A",X"54",X"46",X"84",X"8A",X"3A",X"90",X"01",
		X"0A",X"00",X"08",X"AC",X"00",X"38",X"F0",X"6E",X"A4",X"00",X"68",X"74",X"BE",X"DC",X"88",X"8F",
		X"05",X"00",X"18",X"A9",X"08",X"34",X"FC",X"66",X"8C",X"FA",X"76",X"7A",X"B1",X"CF",X"94",X"92",
		X"07",X"00",X"38",X"BA",X"EC",X"06",X"34",X"0C",X"9C",X"1E",X"76",X"72",X"EF",X"58",X"B3",X"D1",
		X"0E",X"00",X"18",X"BA",X"48",X"06",X"14",X"0C",X"5C",X"1E",X"76",X"72",X"EF",X"58",X"00",X"00",
		X"08",X"00",X"04",X"BA",X"48",X"06",X"14",X"0C",X"5C",X"1E",X"3E",X"72",X"E3",X"58",X"00",X"00",
		X"0A",X"05",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"92",X"54",X"22",X"35",X"00",X"00",
		X"08",X"08",X"00",X"A3",X"E8",X"F0",X"E8",X"08",X"F4",X"F8",X"8E",X"54",X"2A",X"40",X"00",X"00",
		X"0E",X"00",X"14",X"A3",X"48",X"F0",X"08",X"08",X"00",X"F8",X"8E",X"54",X"2A",X"40",X"00",X"00",
		X"01",X"00",X"E0",X"2F",X"00",X"00",X"00",X"00",X"00",X"00",X"4A",X"06",X"62",X"73",X"00",X"00",
		X"03",X"00",X"10",X"6B",X"00",X"00",X"00",X"00",X"00",X"00",X"4A",X"06",X"62",X"73",X"00",X"00",
		X"0C",X"00",X"00",X"00",X"48",X"06",X"00",X"3C",X"40",X"70",X"00",X"6C",X"D6",X"28",X"00",X"00",
		X"0B",X"00",X"40",X"00",X"14",X"20",X"04",X"22",X"D0",X"4A",X"1A",X"5A",X"86",X"F7",X"00",X"00",
		X"01",X"00",X"10",X"FA",X"C4",X"2A",X"34",X"32",X"94",X"34",X"9E",X"0A",X"00",X"E3",X"00",X"00",
		X"08",X"00",X"00",X"FA",X"C4",X"2A",X"34",X"32",X"94",X"34",X"3A",X"0A",X"C0",X"E3",X"00",X"00",
		X"08",X"03",X"00",X"91",X"48",X"7C",X"00",X"58",X"40",X"60",X"F8",X"50",X"C0",X"65",X"00",X"00",
		X"08",X"00",X"00",X"60",X"48",X"7C",X"00",X"58",X"40",X"60",X"F8",X"50",X"C0",X"65",X"00",X"00",
		X"07",X"00",X"18",X"47",X"B0",X"7A",X"F4",X"00",X"98",X"6E",X"CC",X"58",X"D4",X"3B",X"00",X"00",
		X"0C",X"02",X"00",X"73",X"74",X"40",X"08",X"58",X"98",X"6A",X"3A",X"74",X"25",X"16",X"00",X"00",
		X"07",X"00",X"20",X"0D",X"20",X"20",X"20",X"1C",X"84",X"5E",X"8C",X"5C",X"86",X"85",X"00",X"00",
		X"09",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"30",X"33",X"DC",X"4E",X"D0",X"30",X"08",X"5E",X"A8",X"46",X"EF",X"DE",X"00",X"00",
		X"0D",X"00",X"18",X"4F",X"04",X"00",X"A0",X"40",X"F0",X"70",X"52",X"52",X"EF",X"73",X"00",X"00",
		X"37",X"00",X"80",X"3E",X"D8",X"00",X"D8",X"70",X"38",X"00",X"18",X"48",X"54",X"F6",X"24",X"06",
		X"04",X"0E",X"00",X"9D",X"60",X"00",X"30",X"00",X"78",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"01",X"10",X"23",X"29",X"EB",X"09",X"F2",X"4D",X"31",X"44",X"BB",X"61",X"A0",X"BC",X"44",
		X"0D",X"04",X"00",X"9F",X"68",X"40",X"30",X"10",X"C8",X"10",X"9C",X"70",X"04",X"48",X"00",X"00",
		X"0A",X"01",X"80",X"E0",X"60",X"50",X"98",X"40",X"80",X"40",X"00",X"00",X"08",X"E8",X"00",X"00",
		X"01",X"01",X"00",X"A6",X"A8",X"10",X"C8",X"30",X"08",X"60",X"10",X"60",X"30",X"36",X"00",X"00",
		X"06",X"03",X"00",X"42",X"A8",X"10",X"C8",X"30",X"08",X"60",X"10",X"60",X"30",X"36",X"00",X"00",
		X"07",X"01",X"00",X"42",X"A8",X"10",X"C8",X"30",X"08",X"60",X"9C",X"60",X"CC",X"36",X"00",X"00",
		X"04",X"00",X"14",X"CE",X"D8",X"10",X"38",X"30",X"78",X"60",X"9C",X"60",X"CC",X"36",X"00",X"00",
		X"0E",X"00",X"40",X"27",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"18",X"0C",X"80",X"00",X"00",
		X"34",X"00",X"E0",X"6F",X"BC",X"76",X"34",X"40",X"74",X"6C",X"02",X"40",X"28",X"D4",X"00",X"00",
		X"02",X"00",X"40",X"62",X"B8",X"72",X"14",X"44",X"80",X"72",X"14",X"32",X"1B",X"DB",X"00",X"00",
		X"0A",X"02",X"80",X"82",X"08",X"32",X"E0",X"42",X"70",X"5E",X"88",X"7E",X"1E",X"34",X"00",X"00",
		X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0D",X"00",X"07",X"00",X"21",X"18",X"C0",X"0C",X"A5",X"05",X"64",X"9C",X"A5",X"3A",X"C0",X"01",
		X"02",X"00",X"06",X"0C",X"21",X"18",X"C0",X"0C",X"A5",X"05",X"4C",X"AC",X"99",X"30",X"C0",X"01",
		X"02",X"01",X"80",X"33",X"B0",X"40",X"68",X"00",X"08",X"40",X"0C",X"00",X"60",X"66",X"00",X"00",
		X"01",X"00",X"10",X"24",X"83",X"D8",X"5E",X"2F",X"1D",X"19",X"80",X"08",X"3F",X"C4",X"35",X"08",
		X"0C",X"00",X"28",X"24",X"83",X"D8",X"5E",X"2F",X"1D",X"19",X"00",X"08",X"63",X"C4",X"00",X"00",
		X"01",X"03",X"00",X"24",X"83",X"D8",X"5E",X"2F",X"1D",X"19",X"98",X"08",X"FF",X"C4",X"00",X"00",
		X"0A",X"00",X"50",X"CB",X"E3",X"D8",X"6E",X"2F",X"55",X"19",X"98",X"08",X"FF",X"C4",X"00",X"00",
		X"03",X"00",X"20",X"29",X"00",X"30",X"00",X"30",X"48",X"10",X"EC",X"00",X"BC",X"82",X"65",X"78",
		X"04",X"00",X"00",X"00",X"00",X"30",X"00",X"30",X"48",X"10",X"EC",X"00",X"BC",X"82",X"65",X"78",
		X"08",X"08",X"00",X"0F",X"40",X"20",X"08",X"50",X"58",X"30",X"00",X"18",X"C0",X"B0",X"F3",X"66",
		X"0B",X"01",X"40",X"79",X"98",X"20",X"D0",X"50",X"D0",X"30",X"00",X"18",X"C0",X"B0",X"F3",X"66",
		X"02",X"00",X"0C",X"F3",X"20",X"20",X"68",X"50",X"70",X"30",X"00",X"18",X"C0",X"B0",X"F3",X"66",
		X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2E",X"00",X"40",X"DF",X"1C",X"24",X"34",X"5A",X"E4",X"4E",X"98",X"3C",X"49",X"41",X"EF",X"0D",
		X"0F",X"00",X"28",X"CC",X"1C",X"24",X"34",X"5A",X"E4",X"4E",X"98",X"3C",X"49",X"41",X"EF",X"0D",
		X"2A",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"92",X"D0",X"00",X"60",X"00",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"06",X"00",X"2A",X"D0",X"00",X"60",X"00",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"30",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"24",X"25",X"BF",
		X"04",X"00",X"20",X"07",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"F8",X"C0",X"26",X"24",X"BE",
		X"03",X"00",X"14",X"0B",X"00",X"00",X"00",X"F0",X"00",X"10",X"00",X"00",X"C0",X"1E",X"27",X"BB",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"3F",X"00",X"20",X"3A",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"01",X"80",X"AF",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"01",X"40",X"A2",X"20",X"00",X"60",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"18",X"A2",X"20",X"00",X"60",X"00",X"14",X"00",X"1E",X"00",X"00",X"00",X"00",X"00",
		X"09",X"0C",X"00",X"AF",X"20",X"00",X"60",X"00",X"14",X"00",X"3C",X"F8",X"F0",X"0E",X"00",X"00",
		X"06",X"02",X"00",X"03",X"14",X"00",X"B0",X"00",X"F4",X"00",X"3C",X"F8",X"F0",X"0E",X"00",X"00",
		X"08",X"03",X"00",X"F5",X"18",X"6C",X"30",X"44",X"F8",X"06",X"84",X"1E",X"45",X"9B",X"00",X"00",
		X"0E",X"00",X"40",X"B2",X"34",X"6C",X"40",X"44",X"24",X"06",X"84",X"1E",X"45",X"9B",X"00",X"00",
		X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"4F",X"0C",X"06",X"0C",X"FC",X"18",X"06",X"EC",X"FE",X"00",X"02",X"00",X"00",
		X"06",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7C",X"00",X"54",X"00",X"00",X"00",
		X"0B",X"01",X"40",X"79",X"98",X"00",X"D0",X"00",X"D0",X"00",X"7C",X"00",X"54",X"00",X"00",X"00",
		X"02",X"00",X"0C",X"F3",X"20",X"00",X"68",X"00",X"70",X"00",X"7C",X"00",X"54",X"00",X"00",X"00",
		X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"2E",X"00",X"40",X"DF",X"1C",X"24",X"34",X"5A",X"E4",X"4E",X"98",X"3C",X"49",X"41",X"EF",X"0D",
		X"0F",X"00",X"28",X"CC",X"1C",X"24",X"34",X"5A",X"E4",X"4E",X"98",X"3C",X"49",X"41",X"EF",X"0D",
		X"2A",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"92",X"D0",X"00",X"60",X"00",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"06",X"00",X"2A",X"D0",X"00",X"60",X"00",X"D8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"30",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"C4",X"24",X"25",X"BF",
		X"04",X"00",X"20",X"07",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"F8",X"C0",X"26",X"24",X"BE",
		X"03",X"00",X"14",X"0B",X"00",X"00",X"00",X"F0",X"00",X"10",X"00",X"00",X"C0",X"1E",X"27",X"BB",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
