---------------------------------------------------------------------------------
-- sp0256 by Dar (darfpga@aol.fr) (14/04/2018)
-- http://darfpga.blogspot.fr
---------------------------------------------------------------------------------
-- Educational use only
-- Do not redistribute synthetized file with roms
-- Do not redistribute roms whatever the form
-- Use at your own risk
---------------------------------------------------------------------------------
--
-- SP0256-al2 prom decoding scheme and speech synthesis algorithm are from :
--
-- Copyright Joseph Zbiciak, all rights reserved.
-- Copyright tim lindner, all rights reserved.
--
-- See C source code and license in sp0256.c from MAME source
--
-- VHDL code is by Dar.
--
---------------------------------------------------------------------------------
-- Original sp0256 prom is bit compressed. I used sp0256.c from MAME to produce
-- an uncompressed and more easy format to be used in FPGA.
--
-- Original prom is 2K, uncompressed prom is 4k.
--
-- Uncompressed format is :
--
--   64 entries table of 3 bytes/entry : adr_msb, adr_lsb, nb_line (nb parts)
--   (1 entry per allophone)
--
--   Each allophone is made of #nb_line parts
--
--   Each part is described by 16 bytes (one line) : 
--  
--    rpt              : repeat nb 
--    amp_msb, amp_lsb : amplitude
--    per              : periode (number of sample to be produced for each rpt)
--    F0|B0|F1|B1|F2|B2|F3|B3|F4|B4|F5|B5 : filtering coefficients
--
---------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sp0256_al2_decoded is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sp0256_al2_decoded is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
-- adr_msb|adr_lsb|nb_line
X"00",X"0C",X"01", -- #00 : 000-002
X"00",X"0D",X"01", -- #01 : 003-005
X"00",X"0E",X"01", -- #02 : 006-008
X"00",X"0F",X"01", -- #03 : 009-00B
X"00",X"10",X"01", -- #04 : 00C-00E
X"00",X"11",X"0A", -- #05 : 00F-011
X"00",X"1B",X"0A", -- #06 : 012-014
X"00",X"25",X"01", -- #07 : 015-017
X"00",X"26",X"03", -- #08 : 018-01A
X"00",X"29",X"03", -- #09 : 01B-01D
X"00",X"2C",X"03", -- #0A : 01E-020
X"00",X"2F",X"03", -- #0B : 021-023
X"00",X"32",X"01", -- #0C : 024-026
X"00",X"33",X"04", -- #0D : 027-029
X"00",X"37",X"06", -- #0E : 02A-02C
X"00",X"3D",X"01", -- #0F : 02D-02F
X"00",X"3E",X"04", -- #10 : 030-032
X"00",X"42",X"03", -- #11 : 033-035
X"00",X"45",X"02", -- #12 : 036-038
X"00",X"47",X"06", -- #13 : 039-03B
X"00",X"4D",X"08", -- #14 : 03C-03E
X"00",X"55",X"02", -- #15 : 03F-041
X"00",X"57",X"03", -- #16 : 042-044
X"00",X"5A",X"01", -- #17 : 045-047
X"00",X"5B",X"03", -- #18 : 048-04A
X"00",X"5E",X"06", -- #19 : 04B-04D
X"00",X"64",X"01", -- #1A : 04E-050
X"00",X"65",X"03", -- #1B : 051-053
X"00",X"68",X"02", -- #1C : 054-056
X"00",X"6A",X"01", -- #1D : 057-059
X"00",X"6B",X"01", -- #1E : 05A-05C
X"00",X"6C",X"03", -- #1F : 05D-05F
X"00",X"6F",X"05", -- #20 : 060-062
X"00",X"74",X"03", -- #21 : 063-065
X"00",X"77",X"03", -- #22 : 066-068
X"00",X"7A",X"03", -- #23 : 069-06B
X"00",X"7D",X"03", -- #24 : 06C-06E
X"00",X"80",X"04", -- #25 : 06F-071
X"00",X"84",X"02", -- #26 : 072-074
X"00",X"86",X"03", -- #27 : 075-077
X"00",X"89",X"01", -- #28 : 078-07A
X"00",X"8A",X"03", -- #29 : 07B-07D
X"00",X"8D",X"04", -- #2A : 07E-080
X"00",X"91",X"03", -- #2B : 081-083
X"00",X"94",X"04", -- #2C : 084-086
X"00",X"98",X"03", -- #2D : 087-089
X"00",X"9B",X"03", -- #2E : 08A-08C
X"00",X"9E",X"0D", -- #2F : 08D-08F
X"00",X"AB",X"04", -- #30 : 090-092
X"00",X"AF",X"04", -- #31 : 093-095
X"00",X"B3",X"03", -- #32 : 096-098
X"00",X"B6",X"09", -- #33 : 099-09B
X"00",X"BF",X"0A", -- #34 : 09C-09E
X"00",X"C9",X"06", -- #35 : 09F-0A1
X"00",X"CF",X"02", -- #36 : 0A2-0A4
X"00",X"D1",X"01", -- #37 : 0A5-0A7
X"00",X"D2",X"06", -- #38 : 0A8-0AA
X"00",X"D8",X"02", -- #39 : 0AB-0AD
X"00",X"DA",X"09", -- #3A : 0AE-0B0
X"00",X"E3",X"09", -- #3B : 0B1-0B3
X"00",X"EC",X"08", -- #3C : 0B4-0B6
X"00",X"F4",X"03", -- #3D : 0B7-0B9
X"00",X"F7",X"03", -- #3E : 0BA-0BC
X"00",X"FA",X"03", -- #3F : 0BD-0BF
-- rpt|amp_msb mp_lsb|per|F0|B0|F1|B1|F2|B2|F3|B3|F4|B4|F5|B5
X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #00.0 : 0C0-0CF
X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #01.0 : 0D0-0DF
X"07",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #02.0 : 0E0-0EF
X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #03.0 : 0F0-0FF
X"1F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #04.0 : 100-10F
X"03",X"01",X"40",X"5B",X"A0",X"60",X"B8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.0 : 110-11F
X"03",X"00",X"C0",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.1 : 120-12F
X"01",X"00",X"50",X"5B",X"A0",X"60",X"A8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.2 : 130-13F
X"03",X"00",X"80",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.3 : 140-14F
X"01",X"00",X"70",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.4 : 150-15F
X"04",X"00",X"A0",X"5B",X"A0",X"60",X"B8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.5 : 160-16F
X"02",X"01",X"C0",X"5B",X"A8",X"60",X"C0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.6 : 170-17F
X"04",X"02",X"80",X"5B",X"A8",X"60",X"D0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.7 : 180-18F
X"02",X"02",X"80",X"5B",X"A8",X"60",X"E0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.8 : 190-19F
X"09",X"01",X"00",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #05.9 : 1A0-1AF
X"01",X"03",X"00",X"5B",X"B0",X"70",X"C8",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.0 : 1B0-1BF
X"01",X"02",X"80",X"5B",X"C8",X"70",X"B0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.1 : 1C0-1CF
X"02",X"03",X"00",X"5B",X"C8",X"70",X"B0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.2 : 1D0-1DF
X"02",X"02",X"80",X"5B",X"B0",X"70",X"C8",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.3 : 1E0-1EF
X"02",X"02",X"00",X"5B",X"C8",X"70",X"F8",X"70",X"B8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.4 : 1F0-1FF
X"02",X"02",X"80",X"5B",X"B0",X"70",X"D0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.5 : 200-20F
X"03",X"03",X"80",X"5B",X"B0",X"70",X"F8",X"70",X"E0",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.6 : 210-21F
X"01",X"03",X"00",X"5B",X"A8",X"70",X"E0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.7 : 220-22F
X"03",X"02",X"80",X"5B",X"A0",X"70",X"E8",X"70",X"00",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.8 : 230-23F
X"02",X"01",X"00",X"5B",X"A0",X"70",X"F0",X"70",X"00",X"60",X"18",X"50",X"3C",X"44",X"00",X"00", -- #06.9 : 240-24F
X"06",X"06",X"00",X"5B",X"00",X"50",X"28",X"50",X"40",X"50",X"F8",X"10",X"E8",X"58",X"AA",X"64", -- #07.0 : 250-25F
X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #08.0 : 260-26F
X"03",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"40",X"FC",X"04",X"CB",X"68", -- #08.1 : 270-27F
X"05",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"20",X"40",X"C5",X"62", -- #08.2 : 280-28F
X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #09.0 : 290-29F
X"04",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"40",X"F4",X"2C",X"BF",X"3B", -- #09.1 : 2A0-2AF
X"06",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"50",X"F8",X"44",X"CF",X"3A", -- #09.2 : 2B0-2BF
X"04",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"18",X"42",X"FA",X"30", -- #0A.0 : 2C0-2CF
X"04",X"01",X"C0",X"5B",X"18",X"60",X"30",X"50",X"38",X"20",X"00",X"10",X"00",X"60",X"E6",X"38", -- #0A.1 : 2D0-2DF
X"04",X"01",X"40",X"5B",X"18",X"50",X"28",X"40",X"40",X"30",X"FC",X"68",X"E8",X"52",X"DD",X"16", -- #0A.2 : 2E0-2EF
X"07",X"00",X"38",X"5B",X"00",X"30",X"18",X"20",X"38",X"40",X"FC",X"60",X"E0",X"2A",X"A1",X"54", -- #0B.0 : 2F0-2FF
X"03",X"00",X"50",X"5B",X"08",X"30",X"20",X"30",X"20",X"10",X"FC",X"68",X"E8",X"1C",X"A2",X"50", -- #0B.1 : 300-30F
X"09",X"00",X"60",X"5B",X"08",X"30",X"20",X"40",X"20",X"10",X"FC",X"68",X"E0",X"24",X"9B",X"5B", -- #0B.2 : 310-31F
X"05",X"06",X"00",X"5B",X"00",X"50",X"10",X"20",X"30",X"50",X"E8",X"60",X"34",X"1E",X"A0",X"6E", -- #0C.0 : 320-32F
X"05",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #0D.0 : 330-33F
X"03",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"28",X"1C",X"4E",X"F4",X"21", -- #0D.1 : 340-34F
X"04",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"1C",X"44",X"EA",X"53", -- #0D.2 : 350-35F
X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"1C",X"46",X"E7",X"5A", -- #0D.3 : 360-36F
X"05",X"00",X"1C",X"5B",X"98",X"60",X"C0",X"60",X"E0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B", -- #0E.0 : 370-37F
X"03",X"00",X"50",X"5B",X"98",X"60",X"C0",X"60",X"E8",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B", -- #0E.1 : 380-38F
X"01",X"00",X"C0",X"5B",X"98",X"60",X"C0",X"60",X"E8",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B", -- #0E.2 : 390-39F
X"02",X"02",X"80",X"5B",X"A0",X"60",X"C0",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B", -- #0E.3 : 3A0-3AF
X"01",X"01",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B", -- #0E.4 : 3B0-3BF
X"02",X"02",X"00",X"5B",X"A0",X"60",X"B8",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B", -- #0E.5 : 3C0-3CF
X"06",X"06",X"00",X"5B",X"F0",X"50",X"18",X"20",X"28",X"60",X"D0",X"60",X"28",X"18",X"A8",X"61", -- #0F.0 : 3D0-3DF
X"06",X"00",X"A0",X"5B",X"F0",X"50",X"C0",X"30",X"E0",X"20",X"00",X"10",X"20",X"44",X"00",X"00", -- #10.0 : 3E0-3EF
X"05",X"00",X"C0",X"5B",X"F0",X"50",X"C0",X"30",X"E0",X"20",X"00",X"10",X"20",X"44",X"00",X"00", -- #10.1 : 3F0-3FF
X"05",X"00",X"E0",X"5B",X"F0",X"50",X"E0",X"30",X"C8",X"20",X"00",X"10",X"20",X"44",X"00",X"00", -- #10.2 : 400-40F
X"04",X"01",X"40",X"5B",X"F0",X"50",X"E0",X"30",X"C8",X"20",X"00",X"10",X"20",X"44",X"00",X"00", -- #10.3 : 410-41F
X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #11.0 : 420-42F
X"01",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"48",X"10",X"40",X"DF",X"3F", -- #11.1 : 430-43F
X"05",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"28",X"40",X"E8",X"3F", -- #11.2 : 440-44F
X"0C",X"00",X"A0",X"5B",X"08",X"30",X"18",X"30",X"38",X"40",X"EC",X"30",X"D4",X"2E",X"CB",X"20", -- #12.0 : 450-45F
X"03",X"02",X"80",X"5B",X"00",X"60",X"18",X"50",X"38",X"50",X"F4",X"08",X"DC",X"5E",X"A1",X"5C", -- #12.1 : 460-46F
X"03",X"06",X"00",X"5B",X"08",X"00",X"28",X"40",X"38",X"40",X"04",X"60",X"F0",X"66",X"A1",X"5A", -- #13.0 : 470-47F
X"03",X"06",X"00",X"5B",X"28",X"40",X"38",X"40",X"08",X"00",X"04",X"50",X"F4",X"62",X"A4",X"57", -- #13.1 : 480-48F
X"02",X"06",X"00",X"5B",X"08",X"10",X"28",X"50",X"38",X"40",X"04",X"48",X"F4",X"64",X"9A",X"62", -- #13.2 : 490-49F
X"03",X"06",X"00",X"5B",X"08",X"20",X"28",X"50",X"38",X"40",X"04",X"38",X"F8",X"60",X"96",X"66", -- #13.3 : 4A0-4AF
X"04",X"04",X"00",X"5B",X"08",X"30",X"28",X"50",X"38",X"50",X"FC",X"20",X"F8",X"62",X"92",X"6E", -- #13.4 : 4B0-4BF
X"04",X"01",X"40",X"5B",X"08",X"40",X"28",X"40",X"38",X"40",X"F8",X"60",X"F4",X"0C",X"90",X"71", -- #13.5 : 4C0-4CF
X"03",X"03",X"00",X"5B",X"A0",X"70",X"E8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.0 : 4D0-4DF
X"01",X"03",X"00",X"5B",X"A0",X"70",X"F0",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.1 : 4E0-4EF
X"03",X"02",X"80",X"5B",X"A0",X"70",X"F0",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.2 : 4F0-4FF
X"01",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"F8",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.3 : 500-50F
X"05",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.4 : 510-51F
X"01",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.5 : 520-52F
X"06",X"00",X"A0",X"5B",X"90",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.6 : 530-53F
X"02",X"00",X"70",X"5B",X"90",X"70",X"F8",X"60",X"F8",X"20",X"04",X"30",X"28",X"52",X"00",X"00", -- #14.7 : 540-54F
X"03",X"02",X"80",X"5B",X"90",X"70",X"E0",X"70",X"00",X"60",X"10",X"10",X"1C",X"56",X"3A",X"49", -- #15.0 : 550-55F
X"02",X"02",X"00",X"5B",X"98",X"70",X"E0",X"70",X"00",X"60",X"10",X"10",X"1C",X"56",X"3A",X"49", -- #15.1 : 560-56F
X"03",X"05",X"00",X"5B",X"98",X"60",X"F0",X"60",X"D8",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C", -- #16.0 : 570-57F
X"02",X"05",X"00",X"5B",X"D0",X"60",X"F0",X"60",X"A0",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C", -- #16.1 : 580-58F
X"02",X"04",X"00",X"5B",X"F0",X"60",X"C8",X"60",X"A0",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C", -- #16.2 : 590-59F
X"08",X"04",X"00",X"5B",X"20",X"50",X"18",X"20",X"40",X"30",X"F8",X"60",X"C0",X"60",X"B2",X"5A", -- #17.0 : 5A0-5AF
X"03",X"05",X"00",X"5B",X"C8",X"60",X"B8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41", -- #18.0 : 5B0-5BF
X"02",X"05",X"00",X"5B",X"C8",X"60",X"B8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41", -- #18.1 : 5C0-5CF
X"02",X"05",X"00",X"5B",X"B8",X"60",X"C8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41", -- #18.2 : 5D0-5DF
X"03",X"01",X"C0",X"5B",X"10",X"50",X"28",X"40",X"30",X"30",X"08",X"30",X"F0",X"64",X"8E",X"70", -- #19.0 : 5E0-5EF
X"02",X"01",X"80",X"5B",X"10",X"50",X"28",X"50",X"38",X"30",X"04",X"28",X"F4",X"5E",X"8C",X"76", -- #19.1 : 5F0-5FF
X"04",X"02",X"80",X"5B",X"08",X"30",X"28",X"40",X"30",X"20",X"08",X"40",X"F4",X"5C",X"90",X"70", -- #19.2 : 600-60F
X"01",X"04",X"00",X"5B",X"10",X"30",X"20",X"50",X"38",X"40",X"00",X"38",X"F0",X"5A",X"95",X"69", -- #19.3 : 610-61F
X"03",X"07",X"00",X"5B",X"20",X"40",X"28",X"40",X"18",X"10",X"00",X"48",X"F0",X"60",X"98",X"69", -- #19.4 : 620-62F
X"01",X"06",X"00",X"5B",X"18",X"30",X"28",X"40",X"20",X"10",X"00",X"48",X"F0",X"5E",X"9C",X"68", -- #19.5 : 630-63F
X"09",X"03",X"00",X"5B",X"F8",X"40",X"20",X"50",X"30",X"50",X"F0",X"20",X"DC",X"4C",X"AE",X"66", -- #1A.0 : 640-64F
X"06",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"28",X"08",X"4E",X"EB",X"0C", -- #1B.0 : 650-65F
X"06",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"38",X"0C",X"3E",X"F1",X"1A", -- #1B.1 : 660-66F
X"02",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"E8",X"F2",X"03",X"3F", -- #1B.2 : 670-67F
X"03",X"00",X"04",X"5B",X"F8",X"30",X"18",X"40",X"40",X"30",X"E4",X"20",X"18",X"04",X"88",X"76", -- #1C.0 : 680-68F
X"01",X"03",X"00",X"5B",X"20",X"50",X"18",X"10",X"30",X"40",X"F8",X"78",X"E0",X"74",X"98",X"6C", -- #1C.1 : 690-69F
X"14",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"24",X"E5",X"3B", -- #1D.0 : 6A0-6AF
X"08",X"02",X"80",X"5B",X"F8",X"70",X"20",X"50",X"28",X"50",X"C0",X"68",X"18",X"06",X"A4",X"5E", -- #1E.0 : 6B0-6BF
X"08",X"02",X"80",X"5B",X"F0",X"60",X"18",X"60",X"20",X"40",X"D8",X"60",X"20",X"0C",X"9D",X"61", -- #1F.0 : 6C0-6CF
X"04",X"03",X"00",X"5B",X"18",X"50",X"20",X"50",X"38",X"30",X"F0",X"60",X"D0",X"66",X"A6",X"53", -- #1F.1 : 6D0-6DF
X"07",X"02",X"00",X"5B",X"18",X"60",X"28",X"50",X"40",X"40",X"F0",X"60",X"C8",X"62",X"9D",X"61", -- #1F.2 : 6E0-6EF
X"08",X"01",X"C0",X"5B",X"B8",X"60",X"D0",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00", -- #20.0 : 6F0-6FF
X"05",X"01",X"00",X"5B",X"B0",X"60",X"C8",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00", -- #20.1 : 700-70F
X"04",X"00",X"A0",X"5B",X"B0",X"60",X"C0",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00", -- #20.2 : 710-71F
X"04",X"00",X"80",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"50",X"0C",X"20",X"20",X"44",X"00",X"00", -- #20.3 : 720-72F
X"07",X"00",X"28",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"50",X"0C",X"20",X"20",X"44",X"00",X"00", -- #20.4 : 730-73F
X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #21.0 : 740-74F
X"03",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"14",X"32",X"E7",X"23", -- #21.1 : 750-75F
X"03",X"06",X"00",X"5B",X"18",X"50",X"20",X"50",X"40",X"30",X"F8",X"60",X"E4",X"72",X"9D",X"5D", -- #21.2 : 760-76F
X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #22.0 : 770-77F
X"05",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"48",X"F4",X"42",X"EA",X"2A", -- #22.1 : 780-78F
X"03",X"01",X"40",X"5B",X"20",X"30",X"30",X"50",X"18",X"10",X"F8",X"68",X"E8",X"58",X"9C",X"68", -- #22.2 : 790-79F
X"06",X"00",X"20",X"5B",X"08",X"30",X"28",X"50",X"50",X"40",X"F0",X"48",X"C8",X"68",X"A8",X"47", -- #23.0 : 7A0-7AF
X"06",X"00",X"E0",X"5B",X"10",X"40",X"28",X"40",X"50",X"50",X"F0",X"40",X"D0",X"1A",X"DE",X"3A", -- #23.1 : 7B0-7BF
X"02",X"01",X"40",X"5B",X"F0",X"60",X"18",X"40",X"20",X"40",X"D0",X"68",X"2C",X"18",X"C7",X"25", -- #23.2 : 7C0-7CF
X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #24.0 : 7D0-7DF
X"03",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"30",X"FC",X"F0",X"FB",X"41", -- #24.1 : 7E0-7EF
X"03",X"03",X"80",X"5B",X"10",X"40",X"20",X"60",X"38",X"30",X"F8",X"30",X"F4",X"5E",X"A1",X"5C", -- #24.2 : 7F0-7FF
X"06",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"50",X"0C",X"0E",X"FB",X"5C", -- #25.0 : 800-80F
X"03",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"18",X"42",X"FA",X"56", -- #25.1 : 810-81F
X"12",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"18",X"4A",X"FC",X"5B", -- #25.2 : 820-82F
X"04",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"10",X"2E",X"F8",X"4C", -- #25.3 : 830-83F
X"07",X"01",X"40",X"5B",X"C0",X"30",X"E0",X"40",X"F8",X"60",X"14",X"58",X"24",X"48",X"00",X"00", -- #26.0 : 840-84F
X"0B",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"42",X"FE",X"3F", -- #26.1 : 850-85F
X"02",X"00",X"38",X"5B",X"08",X"40",X"20",X"30",X"38",X"30",X"DC",X"48",X"BC",X"58",X"A4",X"54", -- #27.0 : 860-86F
X"03",X"00",X"60",X"5B",X"D0",X"60",X"10",X"70",X"20",X"30",X"BC",X"60",X"1C",X"08",X"A1",X"5D", -- #27.1 : 870-87F
X"04",X"00",X"A0",X"5B",X"D0",X"50",X"10",X"60",X"18",X"50",X"BC",X"60",X"20",X"0E",X"A3",X"5C", -- #27.2 : 880-88F
X"11",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"38",X"04",X"28",X"E3",X"27", -- #28.0 : 890-89F
X"12",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #29.0 : 8A0-8AF
X"01",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"30",X"04",X"12",X"DE",X"56", -- #29.1 : 8B0-8BF
X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"28",X"F4",X"1E",X"DC",X"49", -- #29.2 : 8C0-8CF
X"07",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #2A.0 : 8D0-8DF
X"01",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"0C",X"62",X"E2",X"37", -- #2A.1 : 8E0-8EF
X"01",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"20",X"10",X"36",X"F9",X"44", -- #2A.2 : 8F0-8FF
X"09",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"28",X"0C",X"44",X"E7",X"1B", -- #2A.3 : 900-90F
X"06",X"04",X"00",X"5B",X"20",X"50",X"40",X"60",X"58",X"50",X"00",X"58",X"DC",X"54",X"A7",X"4D", -- #2B.0 : 910-91F
X"09",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"58",X"EC",X"00",X"21",X"30", -- #2B.1 : 920-92F
X"04",X"05",X"00",X"5B",X"20",X"50",X"40",X"50",X"48",X"40",X"00",X"40",X"DC",X"60",X"B9",X"37", -- #2B.2 : 930-93F
X"05",X"03",X"80",X"5B",X"D8",X"40",X"B8",X"40",X"F8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A", -- #2C.0 : 940-94F
X"03",X"02",X"00",X"5B",X"F0",X"40",X"B0",X"40",X"D8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A", -- #2C.1 : 950-95F
X"06",X"01",X"C0",X"5B",X"B0",X"40",X"F0",X"40",X"D8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A", -- #2C.2 : 960-96F
X"08",X"01",X"40",X"5B",X"F0",X"40",X"B0",X"40",X"D0",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A", -- #2C.3 : 970-97F
X"03",X"00",X"C0",X"5B",X"98",X"60",X"C8",X"60",X"08",X"40",X"18",X"30",X"28",X"44",X"2E",X"25", -- #2D.0 : 980-98F
X"03",X"02",X"80",X"5B",X"A0",X"60",X"C8",X"60",X"08",X"40",X"18",X"30",X"28",X"44",X"2E",X"25", -- #2D.1 : 990-99F
X"03",X"02",X"00",X"5B",X"A0",X"60",X"C0",X"60",X"00",X"40",X"18",X"30",X"28",X"44",X"2E",X"25", -- #2D.2 : 9A0-9AF
X"05",X"00",X"28",X"5B",X"F8",X"20",X"18",X"40",X"28",X"30",X"C0",X"38",X"10",X"F8",X"A0",X"5A", -- #2E.0 : 9B0-9BF
X"05",X"00",X"38",X"5B",X"08",X"30",X"20",X"60",X"38",X"40",X"FC",X"08",X"B0",X"50",X"9E",X"5F", -- #2E.1 : 9C0-9CF
X"06",X"00",X"50",X"5B",X"00",X"50",X"18",X"60",X"20",X"50",X"A8",X"70",X"14",X"02",X"93",X"72", -- #2E.2 : 9D0-9DF
X"03",X"02",X"80",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.0 : 9E0-9EF
X"02",X"02",X"80",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.1 : 9F0-9FF
X"02",X"01",X"C0",X"5B",X"A0",X"60",X"E8",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.2 : A00-A0F
X"02",X"02",X"80",X"5B",X"A0",X"60",X"E0",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.3 : A10-A1F
X"02",X"03",X"00",X"5B",X"A8",X"60",X"E0",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.4 : A20-A2F
X"02",X"02",X"80",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.5 : A30-A3F
X"03",X"02",X"00",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.6 : A40-A4F
X"01",X"01",X"C0",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.7 : A50-A5F
X"03",X"00",X"E0",X"5B",X"A8",X"60",X"D0",X"60",X"E0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.8 : A60-A6F
X"01",X"00",X"80",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.9 : A70-A7F
X"02",X"00",X"C0",X"5B",X"A8",X"60",X"D0",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.A : A80-A8F
X"01",X"00",X"70",X"5B",X"A8",X"60",X"D0",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.B : A90-A9F
X"03",X"00",X"50",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59", -- #2F.C : AA0-AAF
X"06",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"FC",X"1C",X"D2",X"28", -- #30.0 : AB0-ABF
X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"38",X"04",X"18",X"B4",X"55", -- #30.1 : AC0-ACF
X"02",X"00",X"C0",X"5B",X"F8",X"40",X"30",X"70",X"20",X"20",X"C4",X"38",X"10",X"FC",X"A3",X"5D", -- #30.2 : AD0-ADF
X"02",X"01",X"40",X"5B",X"F8",X"60",X"28",X"50",X"28",X"50",X"B0",X"68",X"1C",X"06",X"A3",X"58", -- #30.3 : AE0-AEF
X"03",X"01",X"C0",X"5B",X"10",X"50",X"28",X"40",X"30",X"30",X"08",X"30",X"F0",X"64",X"8E",X"70", -- #31.0 : AF0-AFF
X"02",X"01",X"80",X"5B",X"10",X"50",X"28",X"50",X"38",X"30",X"04",X"28",X"F4",X"5E",X"8C",X"76", -- #31.1 : B00-B0F
X"04",X"02",X"80",X"5B",X"08",X"30",X"28",X"40",X"30",X"20",X"08",X"40",X"F4",X"5C",X"90",X"70", -- #31.2 : B10-B1F
X"01",X"04",X"00",X"5B",X"10",X"30",X"20",X"50",X"38",X"40",X"00",X"38",X"F0",X"5A",X"95",X"69", -- #31.3 : B20-B2F
X"05",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #32.0 : B30-B3F
X"05",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"40",X"08",X"4E",X"E4",X"19", -- #32.1 : B40-B4F
X"0D",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"50",X"10",X"66",X"F6",X"49", -- #32.2 : B50-B5F
X"01",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"30",X"20",X"E4",X"60",X"CC",X"68",X"A5",X"5F", -- #33.0 : B60-B6F
X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"28",X"10",X"E4",X"58",X"D0",X"60",X"A5",X"5F", -- #33.1 : B70-B7F
X"01",X"02",X"80",X"5B",X"E0",X"60",X"18",X"40",X"20",X"40",X"D0",X"60",X"24",X"12",X"A8",X"5B", -- #33.2 : B80-B8F
X"01",X"02",X"00",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"20",X"0A",X"A3",X"63", -- #33.3 : B90-B9F
X"01",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D0",X"68",X"20",X"0A",X"A5",X"61", -- #33.4 : BA0-BAF
X"02",X"02",X"00",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"24",X"12",X"A2",X"69", -- #33.5 : BB0-BBF
X"01",X"01",X"40",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D4",X"68",X"1C",X"0A",X"A0",X"6E", -- #33.6 : BC0-BCF
X"02",X"00",X"E0",X"5B",X"18",X"60",X"20",X"20",X"20",X"10",X"E0",X"60",X"D4",X"68",X"A0",X"6E", -- #33.7 : BD0-BDF
X"01",X"01",X"00",X"5B",X"18",X"60",X"18",X"20",X"30",X"20",X"E4",X"60",X"D4",X"6A",X"A3",X"63", -- #33.8 : BE0-BEF
X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"30",X"20",X"E4",X"60",X"CC",X"68",X"A5",X"5F", -- #34.0 : BF0-BFF
X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"28",X"10",X"E4",X"58",X"D0",X"60",X"A5",X"5F", -- #34.1 : C00-C0F
X"02",X"02",X"00",X"5B",X"E0",X"60",X"18",X"40",X"28",X"40",X"D0",X"60",X"24",X"10",X"A9",X"59", -- #34.2 : C10-C1F
X"02",X"02",X"00",X"5B",X"E0",X"60",X"18",X"40",X"20",X"40",X"D0",X"60",X"24",X"12",X"A8",X"5B", -- #34.3 : C20-C2F
X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"20",X"0A",X"A3",X"63", -- #34.4 : C30-C3F
X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D0",X"68",X"20",X"0A",X"A5",X"61", -- #34.5 : C40-C4F
X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"24",X"12",X"A2",X"69", -- #34.6 : C50-C5F
X"03",X"01",X"40",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D4",X"68",X"1C",X"0A",X"A0",X"6E", -- #34.7 : C60-C6F
X"03",X"00",X"C0",X"5B",X"18",X"60",X"20",X"20",X"20",X"10",X"E0",X"60",X"D4",X"68",X"A0",X"6E", -- #34.8 : C70-C7F
X"03",X"00",X"E0",X"5B",X"18",X"60",X"18",X"20",X"30",X"20",X"E4",X"60",X"D4",X"6A",X"A3",X"63", -- #34.9 : C80-C8F
X"03",X"02",X"80",X"5B",X"A8",X"60",X"C0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #35.0 : C90-C9F
X"03",X"02",X"00",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #35.1 : CA0-CAF
X"01",X"01",X"C0",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #35.2 : CB0-CBF
X"05",X"00",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #35.3 : CC0-CCF
X"01",X"00",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #35.4 : CD0-CDF
X"06",X"00",X"70",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00", -- #35.5 : CE0-CEF
X"11",X"00",X"A0",X"5B",X"08",X"30",X"18",X"30",X"38",X"40",X"EC",X"30",X"D4",X"2E",X"CB",X"20", -- #36.0 : CF0-CFF
X"03",X"02",X"80",X"5B",X"00",X"60",X"18",X"50",X"38",X"50",X"F4",X"08",X"DC",X"5E",X"A1",X"5C", -- #36.1 : D00-D0F
X"0A",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"40",X"20",X"38",X"E3",X"29", -- #37.0 : D10-D1F
X"04",X"00",X"A0",X"5B",X"00",X"30",X"18",X"20",X"38",X"40",X"FC",X"60",X"E0",X"2A",X"A1",X"54", -- #38.0 : D20-D2F
X"02",X"00",X"C0",X"5B",X"08",X"30",X"20",X"30",X"20",X"10",X"FC",X"68",X"E8",X"1C",X"A2",X"50", -- #38.1 : D30-D3F
X"02",X"00",X"C0",X"5B",X"08",X"30",X"20",X"40",X"20",X"10",X"FC",X"68",X"E0",X"24",X"9B",X"5B", -- #38.2 : D40-D4F
X"03",X"06",X"00",X"5B",X"10",X"40",X"18",X"40",X"30",X"30",X"F8",X"68",X"DC",X"62",X"A8",X"50", -- #38.3 : D50-D5F
X"01",X"06",X"00",X"5B",X"10",X"20",X"18",X"40",X"30",X"40",X"F8",X"68",X"D4",X"6E",X"AC",X"55", -- #38.4 : D60-D6F
X"03",X"06",X"00",X"5B",X"20",X"50",X"18",X"10",X"30",X"40",X"F8",X"70",X"D0",X"6A",X"AC",X"58", -- #38.5 : D70-D7F
X"0E",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"00",X"1E",X"C1",X"48", -- #39.0 : D80-D8F
X"04",X"00",X"C0",X"5B",X"00",X"40",X"20",X"60",X"38",X"50",X"E8",X"18",X"E0",X"0A",X"C2",X"49", -- #39.1 : D90-D9F
X"02",X"00",X"60",X"5B",X"A0",X"60",X"A8",X"60",X"F8",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.0 : DA0-DAF
X"01",X"00",X"40",X"5B",X"A0",X"60",X"A8",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.1 : DB0-DBF
X"03",X"00",X"50",X"5B",X"A0",X"60",X"A8",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.2 : DC0-DCF
X"03",X"00",X"E0",X"5B",X"A0",X"60",X"B0",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.3 : DD0-DDF
X"05",X"01",X"40",X"5B",X"A0",X"60",X"C0",X"60",X"E8",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.4 : DE0-DEF
X"04",X"01",X"C0",X"5B",X"A8",X"60",X"C8",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.5 : DF0-DFF
X"04",X"01",X"C0",X"5B",X"A8",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.6 : E00-E0F
X"01",X"00",X"E0",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.7 : E10-E1F
X"03",X"00",X"60",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57", -- #3A.8 : E20-E2F
X"02",X"01",X"00",X"5B",X"18",X"60",X"28",X"40",X"10",X"00",X"F0",X"48",X"BC",X"64",X"AC",X"59", -- #3B.0 : E30-E3F
X"02",X"01",X"40",X"5B",X"10",X"60",X"20",X"40",X"18",X"10",X"F0",X"48",X"BC",X"62",X"AF",X"56", -- #3B.1 : E40-E4F
X"02",X"01",X"80",X"5B",X"10",X"50",X"20",X"30",X"20",X"10",X"EC",X"48",X"C0",X"5E",X"B0",X"56", -- #3B.2 : E50-E5F
X"02",X"01",X"40",X"5B",X"F0",X"50",X"10",X"60",X"20",X"50",X"C0",X"60",X"10",X"02",X"B6",X"51", -- #3B.3 : E60-E6F
X"02",X"01",X"40",X"5B",X"E8",X"60",X"18",X"60",X"28",X"50",X"C4",X"60",X"04",X"00",X"B8",X"4A", -- #3B.4 : E70-E7F
X"03",X"01",X"40",X"5B",X"18",X"60",X"10",X"00",X"20",X"30",X"E8",X"58",X"C8",X"62",X"B5",X"54", -- #3B.5 : E80-E8F
X"03",X"00",X"E0",X"5B",X"00",X"00",X"18",X"60",X"30",X"50",X"E4",X"60",X"CC",X"58",X"B5",X"56", -- #3B.6 : E90-E9F
X"03",X"00",X"C0",X"5B",X"00",X"00",X"18",X"60",X"28",X"40",X"E4",X"60",X"D0",X"5C",X"B2",X"59", -- #3B.7 : EA0-EAF
X"03",X"00",X"80",X"5B",X"E8",X"60",X"10",X"60",X"20",X"20",X"CC",X"60",X"04",X"FC",X"B2",X"55", -- #3B.8 : EB0-EBF
X"03",X"03",X"80",X"5B",X"90",X"70",X"F0",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.0 : EC0-ECF
X"02",X"04",X"00",X"5B",X"90",X"70",X"F8",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.1 : ED0-EDF
X"03",X"05",X"00",X"5B",X"90",X"70",X"F8",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.2 : EE0-EEF
X"02",X"02",X"80",X"5B",X"90",X"70",X"F0",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.3 : EF0-EFF
X"03",X"02",X"80",X"5B",X"98",X"70",X"E8",X"50",X"F8",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.4 : F00-F0F
X"04",X"01",X"80",X"5B",X"A0",X"70",X"E0",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.5 : F10-F1F
X"05",X"01",X"80",X"5B",X"A0",X"70",X"D8",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.6 : F20-F2F
X"05",X"01",X"40",X"5B",X"A0",X"70",X"D8",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41", -- #3C.7 : F30-F3F
X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #3D.0 : F40-F4F
X"04",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"E0",X"40",X"E6",X"1C", -- #3D.1 : F50-F5F
X"02",X"01",X"80",X"5B",X"F8",X"40",X"18",X"60",X"38",X"50",X"F8",X"18",X"D8",X"5C",X"A1",X"70", -- #3D.2 : F60-F6F
X"05",X"03",X"00",X"5B",X"18",X"40",X"28",X"50",X"20",X"20",X"FC",X"68",X"C4",X"60",X"A3",X"64", -- #3E.0 : F70-F7F
X"03",X"01",X"80",X"5B",X"10",X"10",X"28",X"60",X"38",X"40",X"FC",X"60",X"C0",X"62",X"A3",X"60", -- #3E.1 : F80-F8F
X"07",X"01",X"00",X"5B",X"28",X"60",X"18",X"10",X"30",X"30",X"00",X"60",X"C0",X"60",X"A0",X"68", -- #3E.2 : F90-F9F
X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", -- #3F.0 : FA0-FAF
X"01",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"FC",X"24",X"DE",X"43", -- #3F.1 : FB0-FBF
X"02",X"05",X"00",X"5B",X"20",X"50",X"30",X"40",X"18",X"10",X"F8",X"68",X"E0",X"6E",X"99",X"6C", -- #3F.2 : FC0-FCF
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --       : FD0-FDF
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00", --       : FE0-FEF
X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00"  --       : FF0-FFF
);
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
