-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb9",
     9 => x"98080b0b",
    10 => x"0bb99c08",
    11 => x"0b0b0bb9",
    12 => x"a0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b9a00c0b",
    16 => x"0b0bb99c",
    17 => x"0c0b0b0b",
    18 => x"b9980c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafe8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b9987080",
    57 => x"c3c8278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e604",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb9a80c",
    65 => x"9f0bb9ac",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b9ac08ff",
    69 => x"05b9ac0c",
    70 => x"b9ac0880",
    71 => x"25eb38b9",
    72 => x"a808ff05",
    73 => x"b9a80cb9",
    74 => x"a8088025",
    75 => x"d738800b",
    76 => x"b9ac0c80",
    77 => x"0bb9a80c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb9a808",
    97 => x"258f3882",
    98 => x"bd2db9a8",
    99 => x"08ff05b9",
   100 => x"a80c82ff",
   101 => x"04b9a808",
   102 => x"b9ac0853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b9a808a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b9ac",
   111 => x"088105b9",
   112 => x"ac0cb9ac",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb9ac0c",
   116 => x"b9a80881",
   117 => x"05b9a80c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b9",
   122 => x"ac088105",
   123 => x"b9ac0cb9",
   124 => x"ac08a02e",
   125 => x"0981068e",
   126 => x"38800bb9",
   127 => x"ac0cb9a8",
   128 => x"088105b9",
   129 => x"a80c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb9b0",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb9b00c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b9",
   169 => x"b0088407",
   170 => x"b9b00c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb594",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b9b00852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b9980c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c8dc12d",
   216 => x"0284050d",
   217 => x"0402fc05",
   218 => x"0dec5192",
   219 => x"710c86a4",
   220 => x"2d82710c",
   221 => x"0284050d",
   222 => x"0402d005",
   223 => x"0d7d5480",
   224 => x"5ba40bec",
   225 => x"0c7352b9",
   226 => x"b451a78e",
   227 => x"2db99808",
   228 => x"7b2e81ab",
   229 => x"38b9b808",
   230 => x"70f80c89",
   231 => x"1580f52d",
   232 => x"8a1680f5",
   233 => x"2d718280",
   234 => x"29058817",
   235 => x"80f52d70",
   236 => x"84808029",
   237 => x"12f40c7e",
   238 => x"ff155c5e",
   239 => x"57555658",
   240 => x"767b2e8b",
   241 => x"38811a77",
   242 => x"812a585a",
   243 => x"76f738f7",
   244 => x"1a5a815b",
   245 => x"80782580",
   246 => x"e6387952",
   247 => x"7651848b",
   248 => x"2dba8052",
   249 => x"b9b451a9",
   250 => x"cd2db998",
   251 => x"08802eb8",
   252 => x"38ba805c",
   253 => x"83fc597b",
   254 => x"7084055d",
   255 => x"087081ff",
   256 => x"0671882a",
   257 => x"7081ff06",
   258 => x"73902a70",
   259 => x"81ff0675",
   260 => x"982ae80c",
   261 => x"e80c58e8",
   262 => x"0c57e80c",
   263 => x"fc1a5a53",
   264 => x"788025d3",
   265 => x"3888af04",
   266 => x"b998085b",
   267 => x"848058b9",
   268 => x"b451a99f",
   269 => x"2dfc8018",
   270 => x"81185858",
   271 => x"87d40486",
   272 => x"b72d800b",
   273 => x"ec0c7a80",
   274 => x"2e8d38b5",
   275 => x"98518fbe",
   276 => x"2d8dc12d",
   277 => x"88dd04b6",
   278 => x"e8518fbe",
   279 => x"2d7ab998",
   280 => x"0c02b005",
   281 => x"0d0402ec",
   282 => x"050d850b",
   283 => x"ec0c8da2",
   284 => x"2d8a8c2d",
   285 => x"81f82d9e",
   286 => x"8d2db998",
   287 => x"08802e80",
   288 => x"f63886f9",
   289 => x"51afe22d",
   290 => x"b598518f",
   291 => x"be2d8dc1",
   292 => x"2d8a982d",
   293 => x"8fce2db5",
   294 => x"c40b80f5",
   295 => x"2d70892b",
   296 => x"9c8006b5",
   297 => x"d00b80f5",
   298 => x"2d70872b",
   299 => x"818006b5",
   300 => x"dc0b80f5",
   301 => x"2d701082",
   302 => x"06747307",
   303 => x"07b5e80b",
   304 => x"80f52d70",
   305 => x"8c2b81e0",
   306 => x"8006b5f4",
   307 => x"0b80f52d",
   308 => x"708f2b82",
   309 => x"80800674",
   310 => x"730707fc",
   311 => x"0c545456",
   312 => x"54525757",
   313 => x"54528652",
   314 => x"b9980885",
   315 => x"38b99808",
   316 => x"5271ec0c",
   317 => x"89910480",
   318 => x"0bb9980c",
   319 => x"0294050d",
   320 => x"0471980c",
   321 => x"04ffb008",
   322 => x"b9980c04",
   323 => x"810bffb0",
   324 => x"0c04800b",
   325 => x"ffb00c04",
   326 => x"02f4050d",
   327 => x"8b9a04b9",
   328 => x"980881f0",
   329 => x"2e098106",
   330 => x"8938810b",
   331 => x"b7cc0c8b",
   332 => x"9a04b998",
   333 => x"0881e02e",
   334 => x"09810689",
   335 => x"38810bb7",
   336 => x"d00c8b9a",
   337 => x"04b99808",
   338 => x"52b7d008",
   339 => x"802e8838",
   340 => x"b9980881",
   341 => x"80055271",
   342 => x"842c728f",
   343 => x"065353b7",
   344 => x"cc08802e",
   345 => x"99387284",
   346 => x"29b78c05",
   347 => x"72138171",
   348 => x"2b700973",
   349 => x"0806730c",
   350 => x"5153538b",
   351 => x"90047284",
   352 => x"29b78c05",
   353 => x"72138371",
   354 => x"2b720807",
   355 => x"720c5353",
   356 => x"800bb7d0",
   357 => x"0c800bb7",
   358 => x"cc0cb9c0",
   359 => x"518c9b2d",
   360 => x"b99808ff",
   361 => x"24fef838",
   362 => x"800bb998",
   363 => x"0c028c05",
   364 => x"0d0402f8",
   365 => x"050db78c",
   366 => x"528f5180",
   367 => x"72708405",
   368 => x"540cff11",
   369 => x"51708025",
   370 => x"f2380288",
   371 => x"050d0402",
   372 => x"f0050d75",
   373 => x"518a922d",
   374 => x"70822cfc",
   375 => x"06b78c11",
   376 => x"72109e06",
   377 => x"71087072",
   378 => x"2a708306",
   379 => x"82742b70",
   380 => x"09740676",
   381 => x"0c545156",
   382 => x"57535153",
   383 => x"8a8c2d71",
   384 => x"b9980c02",
   385 => x"90050d04",
   386 => x"02fc050d",
   387 => x"72518071",
   388 => x"0c800b84",
   389 => x"120c0284",
   390 => x"050d0402",
   391 => x"f0050d75",
   392 => x"70088412",
   393 => x"08535353",
   394 => x"ff547171",
   395 => x"2ea8388a",
   396 => x"922d8413",
   397 => x"08708429",
   398 => x"14881170",
   399 => x"087081ff",
   400 => x"06841808",
   401 => x"81118706",
   402 => x"841a0c53",
   403 => x"51555151",
   404 => x"518a8c2d",
   405 => x"715473b9",
   406 => x"980c0290",
   407 => x"050d0402",
   408 => x"f8050d8a",
   409 => x"922de008",
   410 => x"708b2a70",
   411 => x"81065152",
   412 => x"5270802e",
   413 => x"9d38b9c0",
   414 => x"08708429",
   415 => x"b9c80573",
   416 => x"81ff0671",
   417 => x"0c5151b9",
   418 => x"c0088111",
   419 => x"8706b9c0",
   420 => x"0c51800b",
   421 => x"b9e80c8a",
   422 => x"852d8a8c",
   423 => x"2d028805",
   424 => x"0d0402fc",
   425 => x"050db9c0",
   426 => x"518c882d",
   427 => x"8bb22d8c",
   428 => x"df518a81",
   429 => x"2d028405",
   430 => x"0d04b9ec",
   431 => x"08b9980c",
   432 => x"0402fc05",
   433 => x"0d8dcb04",
   434 => x"8a982d80",
   435 => x"f6518bcf",
   436 => x"2db99808",
   437 => x"f33880da",
   438 => x"518bcf2d",
   439 => x"b99808e8",
   440 => x"38b99808",
   441 => x"b7d80cb9",
   442 => x"98085184",
   443 => x"f02d0284",
   444 => x"050d0402",
   445 => x"ec050d76",
   446 => x"54805287",
   447 => x"0b881580",
   448 => x"f52d5653",
   449 => x"74722483",
   450 => x"38a05372",
   451 => x"5182f92d",
   452 => x"81128b15",
   453 => x"80f52d54",
   454 => x"52727225",
   455 => x"de380294",
   456 => x"050d0402",
   457 => x"f0050db9",
   458 => x"ec085481",
   459 => x"f82d800b",
   460 => x"b9f00c73",
   461 => x"08802e81",
   462 => x"8038820b",
   463 => x"b9ac0cb9",
   464 => x"f0088f06",
   465 => x"b9a80c73",
   466 => x"08527183",
   467 => x"2e963871",
   468 => x"83268938",
   469 => x"71812eaf",
   470 => x"388fa404",
   471 => x"71852e9f",
   472 => x"388fa404",
   473 => x"881480f5",
   474 => x"2d841508",
   475 => x"b3e05354",
   476 => x"5285fe2d",
   477 => x"71842913",
   478 => x"70085252",
   479 => x"8fa80473",
   480 => x"518df32d",
   481 => x"8fa404b7",
   482 => x"d4088815",
   483 => x"082c7081",
   484 => x"06515271",
   485 => x"802e8738",
   486 => x"b3e4518f",
   487 => x"a104b3e8",
   488 => x"5185fe2d",
   489 => x"84140851",
   490 => x"85fe2db9",
   491 => x"f0088105",
   492 => x"b9f00c8c",
   493 => x"14548eb3",
   494 => x"04029005",
   495 => x"0d0471b9",
   496 => x"ec0c8ea3",
   497 => x"2db9f008",
   498 => x"ff05b9f4",
   499 => x"0c0402e8",
   500 => x"050db9ec",
   501 => x"08b9f808",
   502 => x"57558751",
   503 => x"8bcf2db9",
   504 => x"9808812a",
   505 => x"70810651",
   506 => x"5271802e",
   507 => x"a0388ff4",
   508 => x"048a982d",
   509 => x"87518bcf",
   510 => x"2db99808",
   511 => x"f438b7d8",
   512 => x"08813270",
   513 => x"b7d80c70",
   514 => x"525284f0",
   515 => x"2d80fe51",
   516 => x"8bcf2db9",
   517 => x"9808802e",
   518 => x"a638b7d8",
   519 => x"08802e91",
   520 => x"38800bb7",
   521 => x"d80c8051",
   522 => x"84f02d90",
   523 => x"b1048a98",
   524 => x"2d80fe51",
   525 => x"8bcf2db9",
   526 => x"9808f338",
   527 => x"86e52db7",
   528 => x"d8089038",
   529 => x"81fd518b",
   530 => x"cf2d81fa",
   531 => x"518bcf2d",
   532 => x"96840481",
   533 => x"f5518bcf",
   534 => x"2db99808",
   535 => x"812a7081",
   536 => x"06515271",
   537 => x"802eaf38",
   538 => x"b9f40852",
   539 => x"71802e89",
   540 => x"38ff12b9",
   541 => x"f40c9196",
   542 => x"04b9f008",
   543 => x"10b9f008",
   544 => x"05708429",
   545 => x"16515288",
   546 => x"1208802e",
   547 => x"8938ff51",
   548 => x"88120852",
   549 => x"712d81f2",
   550 => x"518bcf2d",
   551 => x"b9980881",
   552 => x"2a708106",
   553 => x"51527180",
   554 => x"2eb138b9",
   555 => x"f008ff11",
   556 => x"b9f40856",
   557 => x"53537372",
   558 => x"25893881",
   559 => x"14b9f40c",
   560 => x"91db0472",
   561 => x"10137084",
   562 => x"29165152",
   563 => x"88120880",
   564 => x"2e8938fe",
   565 => x"51881208",
   566 => x"52712d81",
   567 => x"fd518bcf",
   568 => x"2db99808",
   569 => x"812a7081",
   570 => x"06515271",
   571 => x"802ead38",
   572 => x"b9f40880",
   573 => x"2e893880",
   574 => x"0bb9f40c",
   575 => x"929c04b9",
   576 => x"f00810b9",
   577 => x"f0080570",
   578 => x"84291651",
   579 => x"52881208",
   580 => x"802e8938",
   581 => x"fd518812",
   582 => x"0852712d",
   583 => x"81fa518b",
   584 => x"cf2db998",
   585 => x"08812a70",
   586 => x"81065152",
   587 => x"71802eae",
   588 => x"38b9f008",
   589 => x"ff115452",
   590 => x"b9f40873",
   591 => x"25883872",
   592 => x"b9f40c92",
   593 => x"de047110",
   594 => x"12708429",
   595 => x"16515288",
   596 => x"1208802e",
   597 => x"8938fc51",
   598 => x"88120852",
   599 => x"712db9f4",
   600 => x"08705354",
   601 => x"73802e8a",
   602 => x"388c15ff",
   603 => x"15555592",
   604 => x"e404820b",
   605 => x"b9ac0c71",
   606 => x"8f06b9a8",
   607 => x"0c81eb51",
   608 => x"8bcf2db9",
   609 => x"9808812a",
   610 => x"70810651",
   611 => x"5271802e",
   612 => x"ad387408",
   613 => x"852e0981",
   614 => x"06a43888",
   615 => x"1580f52d",
   616 => x"ff055271",
   617 => x"881681b7",
   618 => x"2d71982b",
   619 => x"52718025",
   620 => x"8838800b",
   621 => x"881681b7",
   622 => x"2d74518d",
   623 => x"f32d81f4",
   624 => x"518bcf2d",
   625 => x"b9980881",
   626 => x"2a708106",
   627 => x"51527180",
   628 => x"2eb33874",
   629 => x"08852e09",
   630 => x"8106aa38",
   631 => x"881580f5",
   632 => x"2d810552",
   633 => x"71881681",
   634 => x"b72d7181",
   635 => x"ff068b16",
   636 => x"80f52d54",
   637 => x"52727227",
   638 => x"87387288",
   639 => x"1681b72d",
   640 => x"74518df3",
   641 => x"2d80da51",
   642 => x"8bcf2db9",
   643 => x"9808812a",
   644 => x"70810651",
   645 => x"5271802e",
   646 => x"81a638b9",
   647 => x"ec08b9f4",
   648 => x"08555373",
   649 => x"802e8a38",
   650 => x"8c13ff15",
   651 => x"555394a3",
   652 => x"04720852",
   653 => x"71822ea6",
   654 => x"38718226",
   655 => x"89387181",
   656 => x"2ea93895",
   657 => x"c0047183",
   658 => x"2eb13871",
   659 => x"842e0981",
   660 => x"0680ed38",
   661 => x"88130851",
   662 => x"8fbe2d95",
   663 => x"c004b9f4",
   664 => x"08518813",
   665 => x"0852712d",
   666 => x"95c00481",
   667 => x"0b881408",
   668 => x"2bb7d408",
   669 => x"32b7d40c",
   670 => x"95960488",
   671 => x"1380f52d",
   672 => x"81058b14",
   673 => x"80f52d53",
   674 => x"54717424",
   675 => x"83388054",
   676 => x"73881481",
   677 => x"b72d8ea3",
   678 => x"2d95c004",
   679 => x"7508802e",
   680 => x"a2387508",
   681 => x"518bcf2d",
   682 => x"b9980881",
   683 => x"06527180",
   684 => x"2e8b38b9",
   685 => x"f4085184",
   686 => x"16085271",
   687 => x"2d881656",
   688 => x"75da3880",
   689 => x"54800bb9",
   690 => x"ac0c738f",
   691 => x"06b9a80c",
   692 => x"a05273b9",
   693 => x"f4082e09",
   694 => x"81069838",
   695 => x"b9f008ff",
   696 => x"05743270",
   697 => x"09810570",
   698 => x"72079f2a",
   699 => x"91713151",
   700 => x"51535371",
   701 => x"5182f92d",
   702 => x"8114548e",
   703 => x"7425c638",
   704 => x"b7d80852",
   705 => x"71b9980c",
   706 => x"0298050d",
   707 => x"0402f405",
   708 => x"0dd45281",
   709 => x"ff720c71",
   710 => x"085381ff",
   711 => x"720c7288",
   712 => x"2b83fe80",
   713 => x"06720870",
   714 => x"81ff0651",
   715 => x"525381ff",
   716 => x"720c7271",
   717 => x"07882b72",
   718 => x"087081ff",
   719 => x"06515253",
   720 => x"81ff720c",
   721 => x"72710788",
   722 => x"2b720870",
   723 => x"81ff0672",
   724 => x"07b9980c",
   725 => x"5253028c",
   726 => x"050d0402",
   727 => x"f4050d74",
   728 => x"767181ff",
   729 => x"06d40c53",
   730 => x"53b9fc08",
   731 => x"85387189",
   732 => x"2b527198",
   733 => x"2ad40c71",
   734 => x"902a7081",
   735 => x"ff06d40c",
   736 => x"5171882a",
   737 => x"7081ff06",
   738 => x"d40c5171",
   739 => x"81ff06d4",
   740 => x"0c72902a",
   741 => x"7081ff06",
   742 => x"d40c51d4",
   743 => x"087081ff",
   744 => x"06515182",
   745 => x"b8bf5270",
   746 => x"81ff2e09",
   747 => x"81069438",
   748 => x"81ff0bd4",
   749 => x"0cd40870",
   750 => x"81ff06ff",
   751 => x"14545151",
   752 => x"71e53870",
   753 => x"b9980c02",
   754 => x"8c050d04",
   755 => x"02fc050d",
   756 => x"81c75181",
   757 => x"ff0bd40c",
   758 => x"ff115170",
   759 => x"8025f438",
   760 => x"0284050d",
   761 => x"0402f405",
   762 => x"0d81ff0b",
   763 => x"d40c9353",
   764 => x"805287fc",
   765 => x"80c15196",
   766 => x"db2db998",
   767 => x"088b3881",
   768 => x"ff0bd40c",
   769 => x"81539892",
   770 => x"0497cc2d",
   771 => x"ff135372",
   772 => x"df3872b9",
   773 => x"980c028c",
   774 => x"050d0402",
   775 => x"ec050d81",
   776 => x"0bb9fc0c",
   777 => x"8454d008",
   778 => x"708f2a70",
   779 => x"81065151",
   780 => x"5372f338",
   781 => x"72d00c97",
   782 => x"cc2db3ec",
   783 => x"5185fe2d",
   784 => x"d008708f",
   785 => x"2a708106",
   786 => x"51515372",
   787 => x"f338810b",
   788 => x"d00cb153",
   789 => x"805284d4",
   790 => x"80c05196",
   791 => x"db2db998",
   792 => x"08812e93",
   793 => x"3872822e",
   794 => x"bd38ff13",
   795 => x"5372e538",
   796 => x"ff145473",
   797 => x"ffb03897",
   798 => x"cc2d83aa",
   799 => x"52849c80",
   800 => x"c85196db",
   801 => x"2db99808",
   802 => x"812e0981",
   803 => x"06923896",
   804 => x"8d2db998",
   805 => x"0883ffff",
   806 => x"06537283",
   807 => x"aa2e9d38",
   808 => x"97e52d99",
   809 => x"b704b3f8",
   810 => x"5185fe2d",
   811 => x"80539b85",
   812 => x"04b49051",
   813 => x"85fe2d80",
   814 => x"549ad704",
   815 => x"81ff0bd4",
   816 => x"0cb15497",
   817 => x"cc2d8fcf",
   818 => x"53805287",
   819 => x"fc80f751",
   820 => x"96db2db9",
   821 => x"980855b9",
   822 => x"9808812e",
   823 => x"0981069b",
   824 => x"3881ff0b",
   825 => x"d40c820a",
   826 => x"52849c80",
   827 => x"e95196db",
   828 => x"2db99808",
   829 => x"802e8d38",
   830 => x"97cc2dff",
   831 => x"135372c9",
   832 => x"389aca04",
   833 => x"81ff0bd4",
   834 => x"0cb99808",
   835 => x"5287fc80",
   836 => x"fa5196db",
   837 => x"2db99808",
   838 => x"b13881ff",
   839 => x"0bd40cd4",
   840 => x"085381ff",
   841 => x"0bd40c81",
   842 => x"ff0bd40c",
   843 => x"81ff0bd4",
   844 => x"0c81ff0b",
   845 => x"d40c7286",
   846 => x"2a708106",
   847 => x"76565153",
   848 => x"729538b9",
   849 => x"9808549a",
   850 => x"d7047382",
   851 => x"2efee238",
   852 => x"ff145473",
   853 => x"feed3873",
   854 => x"b9fc0c73",
   855 => x"8b388152",
   856 => x"87fc80d0",
   857 => x"5196db2d",
   858 => x"81ff0bd4",
   859 => x"0cd00870",
   860 => x"8f2a7081",
   861 => x"06515153",
   862 => x"72f33872",
   863 => x"d00c81ff",
   864 => x"0bd40c81",
   865 => x"5372b998",
   866 => x"0c029405",
   867 => x"0d0402e8",
   868 => x"050d7855",
   869 => x"805681ff",
   870 => x"0bd40cd0",
   871 => x"08708f2a",
   872 => x"70810651",
   873 => x"515372f3",
   874 => x"3882810b",
   875 => x"d00c81ff",
   876 => x"0bd40c77",
   877 => x"5287fc80",
   878 => x"d15196db",
   879 => x"2d80dbc6",
   880 => x"df54b998",
   881 => x"08802e8a",
   882 => x"38b4b051",
   883 => x"85fe2d9c",
   884 => x"a50481ff",
   885 => x"0bd40cd4",
   886 => x"087081ff",
   887 => x"06515372",
   888 => x"81fe2e09",
   889 => x"81069d38",
   890 => x"80ff5396",
   891 => x"8d2db998",
   892 => x"08757084",
   893 => x"05570cff",
   894 => x"13537280",
   895 => x"25ed3881",
   896 => x"569c8a04",
   897 => x"ff145473",
   898 => x"c93881ff",
   899 => x"0bd40c81",
   900 => x"ff0bd40c",
   901 => x"d008708f",
   902 => x"2a708106",
   903 => x"51515372",
   904 => x"f33872d0",
   905 => x"0c75b998",
   906 => x"0c029805",
   907 => x"0d0402e8",
   908 => x"050d7779",
   909 => x"7b585555",
   910 => x"80537276",
   911 => x"25a33874",
   912 => x"70810556",
   913 => x"80f52d74",
   914 => x"70810556",
   915 => x"80f52d52",
   916 => x"5271712e",
   917 => x"86388151",
   918 => x"9ce30481",
   919 => x"13539cba",
   920 => x"04805170",
   921 => x"b9980c02",
   922 => x"98050d04",
   923 => x"02ec050d",
   924 => x"76557480",
   925 => x"2ebe389a",
   926 => x"1580e02d",
   927 => x"51aaa62d",
   928 => x"b99808b9",
   929 => x"980880c0",
   930 => x"b00cb998",
   931 => x"08545480",
   932 => x"c08c0880",
   933 => x"2e993894",
   934 => x"1580e02d",
   935 => x"51aaa62d",
   936 => x"b9980890",
   937 => x"2b83fff0",
   938 => x"0a067075",
   939 => x"07515372",
   940 => x"80c0b00c",
   941 => x"80c0b008",
   942 => x"5372802e",
   943 => x"9d3880c0",
   944 => x"8408fe14",
   945 => x"712980c0",
   946 => x"98080580",
   947 => x"c0b40c70",
   948 => x"842b80c0",
   949 => x"900c549e",
   950 => x"880480c0",
   951 => x"9c0880c0",
   952 => x"b00c80c0",
   953 => x"a00880c0",
   954 => x"b40c80c0",
   955 => x"8c08802e",
   956 => x"8b3880c0",
   957 => x"8408842b",
   958 => x"539e8304",
   959 => x"80c0a408",
   960 => x"842b5372",
   961 => x"80c0900c",
   962 => x"0294050d",
   963 => x"0402d805",
   964 => x"0d800b80",
   965 => x"c08c0c84",
   966 => x"54989b2d",
   967 => x"b9980880",
   968 => x"2e9538ba",
   969 => x"80528051",
   970 => x"9b8e2db9",
   971 => x"9808802e",
   972 => x"8638fe54",
   973 => x"9ebf04ff",
   974 => x"14547380",
   975 => x"24db3873",
   976 => x"8c38b4c0",
   977 => x"5185fe2d",
   978 => x"7355a3e1",
   979 => x"04805681",
   980 => x"0b80c0b8",
   981 => x"0c8853b4",
   982 => x"d452bab6",
   983 => x"519cae2d",
   984 => x"b9980876",
   985 => x"2e098106",
   986 => x"8838b998",
   987 => x"0880c0b8",
   988 => x"0c8853b4",
   989 => x"e052bad2",
   990 => x"519cae2d",
   991 => x"b9980888",
   992 => x"38b99808",
   993 => x"80c0b80c",
   994 => x"80c0b808",
   995 => x"802e80f6",
   996 => x"38bdc60b",
   997 => x"80f52dbd",
   998 => x"c70b80f5",
   999 => x"2d71982b",
  1000 => x"71902b07",
  1001 => x"bdc80b80",
  1002 => x"f52d7088",
  1003 => x"2b7207bd",
  1004 => x"c90b80f5",
  1005 => x"2d7107bd",
  1006 => x"fe0b80f5",
  1007 => x"2dbdff0b",
  1008 => x"80f52d71",
  1009 => x"882b0753",
  1010 => x"5f54525a",
  1011 => x"56575573",
  1012 => x"81abaa2e",
  1013 => x"0981068d",
  1014 => x"387551a9",
  1015 => x"f62db998",
  1016 => x"08569ff2",
  1017 => x"047382d4",
  1018 => x"d52e8738",
  1019 => x"b4ec51a0",
  1020 => x"b404ba80",
  1021 => x"5275519b",
  1022 => x"8e2db998",
  1023 => x"0855b998",
  1024 => x"08802e83",
  1025 => x"dc388853",
  1026 => x"b4e052ba",
  1027 => x"d2519cae",
  1028 => x"2db99808",
  1029 => x"8a38810b",
  1030 => x"80c08c0c",
  1031 => x"a0ba0488",
  1032 => x"53b4d452",
  1033 => x"bab6519c",
  1034 => x"ae2db998",
  1035 => x"08802e8a",
  1036 => x"38b58051",
  1037 => x"85fe2da1",
  1038 => x"9404bdfe",
  1039 => x"0b80f52d",
  1040 => x"547380d5",
  1041 => x"2e098106",
  1042 => x"80ca38bd",
  1043 => x"ff0b80f5",
  1044 => x"2d547381",
  1045 => x"aa2e0981",
  1046 => x"06ba3880",
  1047 => x"0bba800b",
  1048 => x"80f52d56",
  1049 => x"547481e9",
  1050 => x"2e833881",
  1051 => x"547481eb",
  1052 => x"2e8c3880",
  1053 => x"5573752e",
  1054 => x"09810682",
  1055 => x"e438ba8b",
  1056 => x"0b80f52d",
  1057 => x"55748d38",
  1058 => x"ba8c0b80",
  1059 => x"f52d5473",
  1060 => x"822e8638",
  1061 => x"8055a3e1",
  1062 => x"04ba8d0b",
  1063 => x"80f52d70",
  1064 => x"80c0840c",
  1065 => x"ff0580c0",
  1066 => x"880cba8e",
  1067 => x"0b80f52d",
  1068 => x"ba8f0b80",
  1069 => x"f52d5876",
  1070 => x"05778280",
  1071 => x"29057080",
  1072 => x"c0940cba",
  1073 => x"900b80f5",
  1074 => x"2d7080c0",
  1075 => x"a80c80c0",
  1076 => x"8c085957",
  1077 => x"5876802e",
  1078 => x"81ac3888",
  1079 => x"53b4e052",
  1080 => x"bad2519c",
  1081 => x"ae2db998",
  1082 => x"0881f638",
  1083 => x"80c08408",
  1084 => x"70842b80",
  1085 => x"c0900c70",
  1086 => x"80c0a40c",
  1087 => x"baa50b80",
  1088 => x"f52dbaa4",
  1089 => x"0b80f52d",
  1090 => x"71828029",
  1091 => x"05baa60b",
  1092 => x"80f52d70",
  1093 => x"84808029",
  1094 => x"12baa70b",
  1095 => x"80f52d70",
  1096 => x"81800a29",
  1097 => x"127080c0",
  1098 => x"ac0c80c0",
  1099 => x"a8087129",
  1100 => x"80c09408",
  1101 => x"057080c0",
  1102 => x"980cbaad",
  1103 => x"0b80f52d",
  1104 => x"baac0b80",
  1105 => x"f52d7182",
  1106 => x"802905ba",
  1107 => x"ae0b80f5",
  1108 => x"2d708480",
  1109 => x"802912ba",
  1110 => x"af0b80f5",
  1111 => x"2d70982b",
  1112 => x"81f00a06",
  1113 => x"72057080",
  1114 => x"c09c0cfe",
  1115 => x"117e2977",
  1116 => x"0580c0a0",
  1117 => x"0c525952",
  1118 => x"43545e51",
  1119 => x"5259525d",
  1120 => x"575957a3",
  1121 => x"da04ba92",
  1122 => x"0b80f52d",
  1123 => x"ba910b80",
  1124 => x"f52d7182",
  1125 => x"80290570",
  1126 => x"80c0900c",
  1127 => x"70a02983",
  1128 => x"ff057089",
  1129 => x"2a7080c0",
  1130 => x"a40cba97",
  1131 => x"0b80f52d",
  1132 => x"ba960b80",
  1133 => x"f52d7182",
  1134 => x"80290570",
  1135 => x"80c0ac0c",
  1136 => x"7b71291e",
  1137 => x"7080c0a0",
  1138 => x"0c7d80c0",
  1139 => x"9c0c7305",
  1140 => x"80c0980c",
  1141 => x"555e5151",
  1142 => x"55558051",
  1143 => x"9cec2d81",
  1144 => x"5574b998",
  1145 => x"0c02a805",
  1146 => x"0d0402ec",
  1147 => x"050d7670",
  1148 => x"872c7180",
  1149 => x"ff065556",
  1150 => x"5480c08c",
  1151 => x"088a3873",
  1152 => x"882c7481",
  1153 => x"ff065455",
  1154 => x"ba805280",
  1155 => x"c0940815",
  1156 => x"519b8e2d",
  1157 => x"b9980854",
  1158 => x"b9980880",
  1159 => x"2eb43880",
  1160 => x"c08c0880",
  1161 => x"2e983872",
  1162 => x"8429ba80",
  1163 => x"05700852",
  1164 => x"53a9f62d",
  1165 => x"b99808f0",
  1166 => x"0a0653a4",
  1167 => x"d0047210",
  1168 => x"ba800570",
  1169 => x"80e02d52",
  1170 => x"53aaa62d",
  1171 => x"b9980853",
  1172 => x"725473b9",
  1173 => x"980c0294",
  1174 => x"050d0402",
  1175 => x"e0050d79",
  1176 => x"70842c80",
  1177 => x"c0b40805",
  1178 => x"718f0652",
  1179 => x"55537289",
  1180 => x"38ba8052",
  1181 => x"73519b8e",
  1182 => x"2d72a029",
  1183 => x"ba800554",
  1184 => x"807480f5",
  1185 => x"2d565374",
  1186 => x"732e8338",
  1187 => x"81537481",
  1188 => x"e52e81ef",
  1189 => x"38817074",
  1190 => x"06545872",
  1191 => x"802e81e3",
  1192 => x"388b1480",
  1193 => x"f52d7083",
  1194 => x"2a790658",
  1195 => x"56769838",
  1196 => x"b7dc0853",
  1197 => x"72883872",
  1198 => x"be800b81",
  1199 => x"b72d76b7",
  1200 => x"dc0c7353",
  1201 => x"a7850475",
  1202 => x"8f2e0981",
  1203 => x"0681b438",
  1204 => x"749f068d",
  1205 => x"29bdf311",
  1206 => x"51538114",
  1207 => x"80f52d73",
  1208 => x"70810555",
  1209 => x"81b72d83",
  1210 => x"1480f52d",
  1211 => x"73708105",
  1212 => x"5581b72d",
  1213 => x"851480f5",
  1214 => x"2d737081",
  1215 => x"055581b7",
  1216 => x"2d871480",
  1217 => x"f52d7370",
  1218 => x"81055581",
  1219 => x"b72d8914",
  1220 => x"80f52d73",
  1221 => x"70810555",
  1222 => x"81b72d8e",
  1223 => x"1480f52d",
  1224 => x"73708105",
  1225 => x"5581b72d",
  1226 => x"901480f5",
  1227 => x"2d737081",
  1228 => x"055581b7",
  1229 => x"2d921480",
  1230 => x"f52d7370",
  1231 => x"81055581",
  1232 => x"b72d9414",
  1233 => x"80f52d73",
  1234 => x"70810555",
  1235 => x"81b72d96",
  1236 => x"1480f52d",
  1237 => x"73708105",
  1238 => x"5581b72d",
  1239 => x"981480f5",
  1240 => x"2d737081",
  1241 => x"055581b7",
  1242 => x"2d9c1480",
  1243 => x"f52d7370",
  1244 => x"81055581",
  1245 => x"b72d9e14",
  1246 => x"80f52d73",
  1247 => x"81b72d77",
  1248 => x"b7dc0c80",
  1249 => x"5372b998",
  1250 => x"0c02a005",
  1251 => x"0d0402cc",
  1252 => x"050d7e60",
  1253 => x"5e5a800b",
  1254 => x"80c0b008",
  1255 => x"80c0b408",
  1256 => x"595c5680",
  1257 => x"5880c090",
  1258 => x"08782e81",
  1259 => x"b038778f",
  1260 => x"06a01757",
  1261 => x"54738f38",
  1262 => x"ba805276",
  1263 => x"51811757",
  1264 => x"9b8e2dba",
  1265 => x"80568076",
  1266 => x"80f52d56",
  1267 => x"5474742e",
  1268 => x"83388154",
  1269 => x"7481e52e",
  1270 => x"80f73881",
  1271 => x"70750655",
  1272 => x"5c73802e",
  1273 => x"80eb388b",
  1274 => x"1680f52d",
  1275 => x"98065978",
  1276 => x"80df388b",
  1277 => x"537c5275",
  1278 => x"519cae2d",
  1279 => x"b9980880",
  1280 => x"d0389c16",
  1281 => x"0851a9f6",
  1282 => x"2db99808",
  1283 => x"841b0c9a",
  1284 => x"1680e02d",
  1285 => x"51aaa62d",
  1286 => x"b99808b9",
  1287 => x"9808881c",
  1288 => x"0cb99808",
  1289 => x"555580c0",
  1290 => x"8c08802e",
  1291 => x"98389416",
  1292 => x"80e02d51",
  1293 => x"aaa62db9",
  1294 => x"9808902b",
  1295 => x"83fff00a",
  1296 => x"06701651",
  1297 => x"5473881b",
  1298 => x"0c787a0c",
  1299 => x"7b54a996",
  1300 => x"04811858",
  1301 => x"80c09008",
  1302 => x"7826fed2",
  1303 => x"3880c08c",
  1304 => x"08802eb0",
  1305 => x"387a51a3",
  1306 => x"ea2db998",
  1307 => x"08b99808",
  1308 => x"80ffffff",
  1309 => x"f806555b",
  1310 => x"7380ffff",
  1311 => x"fff82e94",
  1312 => x"38b99808",
  1313 => x"fe0580c0",
  1314 => x"84082980",
  1315 => x"c0980805",
  1316 => x"57a7a304",
  1317 => x"805473b9",
  1318 => x"980c02b4",
  1319 => x"050d0402",
  1320 => x"f4050d74",
  1321 => x"70088105",
  1322 => x"710c7008",
  1323 => x"80c08808",
  1324 => x"06535371",
  1325 => x"8e388813",
  1326 => x"0851a3ea",
  1327 => x"2db99808",
  1328 => x"88140c81",
  1329 => x"0bb9980c",
  1330 => x"028c050d",
  1331 => x"0402f005",
  1332 => x"0d758811",
  1333 => x"08fe0580",
  1334 => x"c0840829",
  1335 => x"80c09808",
  1336 => x"11720880",
  1337 => x"c0880806",
  1338 => x"05795553",
  1339 => x"54549b8e",
  1340 => x"2d029005",
  1341 => x"0d0402f4",
  1342 => x"050d7470",
  1343 => x"882a83fe",
  1344 => x"80067072",
  1345 => x"982a0772",
  1346 => x"882b87fc",
  1347 => x"80800673",
  1348 => x"982b81f0",
  1349 => x"0a067173",
  1350 => x"0707b998",
  1351 => x"0c565153",
  1352 => x"51028c05",
  1353 => x"0d0402f8",
  1354 => x"050d028e",
  1355 => x"0580f52d",
  1356 => x"74882b07",
  1357 => x"7083ffff",
  1358 => x"06b9980c",
  1359 => x"51028805",
  1360 => x"0d0402f4",
  1361 => x"050d7476",
  1362 => x"78535452",
  1363 => x"80712597",
  1364 => x"38727081",
  1365 => x"055480f5",
  1366 => x"2d727081",
  1367 => x"055481b7",
  1368 => x"2dff1151",
  1369 => x"70eb3880",
  1370 => x"7281b72d",
  1371 => x"028c050d",
  1372 => x"0402e805",
  1373 => x"0d775680",
  1374 => x"70565473",
  1375 => x"7624b338",
  1376 => x"80c09008",
  1377 => x"742eab38",
  1378 => x"7351a4db",
  1379 => x"2db99808",
  1380 => x"b9980809",
  1381 => x"810570b9",
  1382 => x"9808079f",
  1383 => x"2a770581",
  1384 => x"17575753",
  1385 => x"53747624",
  1386 => x"893880c0",
  1387 => x"90087426",
  1388 => x"d73872b9",
  1389 => x"980c0298",
  1390 => x"050d0402",
  1391 => x"f0050db9",
  1392 => x"94081651",
  1393 => x"aaf12db9",
  1394 => x"9808802e",
  1395 => x"9c388b53",
  1396 => x"b9980852",
  1397 => x"be8051aa",
  1398 => x"c22d80c0",
  1399 => x"bc085473",
  1400 => x"802e8638",
  1401 => x"be805173",
  1402 => x"2d029005",
  1403 => x"0d0402dc",
  1404 => x"050d8070",
  1405 => x"5a5574b9",
  1406 => x"940825b1",
  1407 => x"3880c090",
  1408 => x"08752ea9",
  1409 => x"387851a4",
  1410 => x"db2db998",
  1411 => x"08098105",
  1412 => x"70b99808",
  1413 => x"079f2a76",
  1414 => x"05811b5b",
  1415 => x"565474b9",
  1416 => x"94082589",
  1417 => x"3880c090",
  1418 => x"087926d9",
  1419 => x"38805578",
  1420 => x"80c09008",
  1421 => x"2781d138",
  1422 => x"7851a4db",
  1423 => x"2db99808",
  1424 => x"802e81a5",
  1425 => x"38b99808",
  1426 => x"8b0580f5",
  1427 => x"2d70842a",
  1428 => x"70810677",
  1429 => x"1078842b",
  1430 => x"be800b80",
  1431 => x"f52d5c5c",
  1432 => x"53515556",
  1433 => x"73802e80",
  1434 => x"c8387416",
  1435 => x"822baeac",
  1436 => x"0bb7e812",
  1437 => x"0c547775",
  1438 => x"311080c0",
  1439 => x"c0115556",
  1440 => x"90747081",
  1441 => x"055681b7",
  1442 => x"2da07481",
  1443 => x"b72d7681",
  1444 => x"ff068116",
  1445 => x"58547380",
  1446 => x"2e89389c",
  1447 => x"53be8052",
  1448 => x"ada9048b",
  1449 => x"53b99808",
  1450 => x"5280c0c2",
  1451 => x"1651ade1",
  1452 => x"04741682",
  1453 => x"2babbb0b",
  1454 => x"b7e8120c",
  1455 => x"547681ff",
  1456 => x"06811658",
  1457 => x"5473802e",
  1458 => x"89389c53",
  1459 => x"be8052ad",
  1460 => x"d8048b53",
  1461 => x"b9980852",
  1462 => x"77753110",
  1463 => x"80c0c005",
  1464 => x"517655aa",
  1465 => x"c22dadfd",
  1466 => x"04749029",
  1467 => x"75317010",
  1468 => x"80c0c005",
  1469 => x"5154b998",
  1470 => x"087481b7",
  1471 => x"2d811959",
  1472 => x"748b24a3",
  1473 => x"38acaf04",
  1474 => x"74902975",
  1475 => x"31701080",
  1476 => x"c0c0058c",
  1477 => x"77315751",
  1478 => x"54807481",
  1479 => x"b72d9e14",
  1480 => x"ff165654",
  1481 => x"74f33802",
  1482 => x"a4050d04",
  1483 => x"02fc050d",
  1484 => x"b9940813",
  1485 => x"51aaf12d",
  1486 => x"b9980880",
  1487 => x"2e8838b9",
  1488 => x"9808519c",
  1489 => x"ec2d800b",
  1490 => x"b9940cab",
  1491 => x"ee2d8ea3",
  1492 => x"2d028405",
  1493 => x"0d0402fc",
  1494 => x"050d7251",
  1495 => x"70fd2ead",
  1496 => x"3870fd24",
  1497 => x"8a3870fc",
  1498 => x"2e80c438",
  1499 => x"afb70470",
  1500 => x"fe2eb138",
  1501 => x"70ff2e09",
  1502 => x"8106bc38",
  1503 => x"b9940851",
  1504 => x"70802eb3",
  1505 => x"38ff11b9",
  1506 => x"940cafb7",
  1507 => x"04b99408",
  1508 => x"f00570b9",
  1509 => x"940c5170",
  1510 => x"80259c38",
  1511 => x"800bb994",
  1512 => x"0cafb704",
  1513 => x"b9940881",
  1514 => x"05b9940c",
  1515 => x"afb704b9",
  1516 => x"94089005",
  1517 => x"b9940cab",
  1518 => x"ee2d8ea3",
  1519 => x"2d028405",
  1520 => x"0d0402fc",
  1521 => x"050d800b",
  1522 => x"b9940cab",
  1523 => x"ee2d8dba",
  1524 => x"2db99808",
  1525 => x"b9840cb7",
  1526 => x"e0518fbe",
  1527 => x"2d028405",
  1528 => x"0d047180",
  1529 => x"c0bc0c04",
  1530 => x"00ffffff",
  1531 => x"ff00ffff",
  1532 => x"ffff00ff",
  1533 => x"ffffff00",
  1534 => x"20203d56",
  1535 => x"6964656f",
  1536 => x"7061632f",
  1537 => x"4f646479",
  1538 => x"73657932",
  1539 => x"3d202000",
  1540 => x"20202020",
  1541 => x"20202020",
  1542 => x"20202020",
  1543 => x"20202020",
  1544 => x"20202020",
  1545 => x"20202000",
  1546 => x"52657365",
  1547 => x"74000000",
  1548 => x"43617267",
  1549 => x"61722043",
  1550 => x"61727475",
  1551 => x"63686f2f",
  1552 => x"466f6e74",
  1553 => x"20100000",
  1554 => x"45786974",
  1555 => x"00000000",
  1556 => x"53797374",
  1557 => x"656d3a20",
  1558 => x"4f647973",
  1559 => x"73657932",
  1560 => x"00000000",
  1561 => x"53797374",
  1562 => x"656d3a20",
  1563 => x"56696465",
  1564 => x"6f706163",
  1565 => x"00000000",
  1566 => x"47373230",
  1567 => x"30204d6f",
  1568 => x"64653a20",
  1569 => x"4f666600",
  1570 => x"47373230",
  1571 => x"30204d6f",
  1572 => x"64653a20",
  1573 => x"436f6e74",
  1574 => x"72617374",
  1575 => x"20310000",
  1576 => x"47373230",
  1577 => x"30204d6f",
  1578 => x"64653a20",
  1579 => x"436f6e74",
  1580 => x"72617374",
  1581 => x"20320000",
  1582 => x"47373230",
  1583 => x"30204d6f",
  1584 => x"64653a20",
  1585 => x"436f6e74",
  1586 => x"72617374",
  1587 => x"20330000",
  1588 => x"47373230",
  1589 => x"30204d6f",
  1590 => x"64653a20",
  1591 => x"436f6e74",
  1592 => x"72617374",
  1593 => x"20340000",
  1594 => x"47373230",
  1595 => x"30204d6f",
  1596 => x"64653a20",
  1597 => x"436f6e74",
  1598 => x"72617374",
  1599 => x"20350000",
  1600 => x"47373230",
  1601 => x"30204d6f",
  1602 => x"64653a20",
  1603 => x"436f6e74",
  1604 => x"72617374",
  1605 => x"20360000",
  1606 => x"47373230",
  1607 => x"30204d6f",
  1608 => x"64653a20",
  1609 => x"436f6e74",
  1610 => x"72617374",
  1611 => x"20370000",
  1612 => x"54686520",
  1613 => x"566f6963",
  1614 => x"653a204f",
  1615 => x"66660000",
  1616 => x"54686520",
  1617 => x"566f6963",
  1618 => x"653a204f",
  1619 => x"6e000000",
  1620 => x"53776170",
  1621 => x"204a6f79",
  1622 => x"3a204f66",
  1623 => x"66000000",
  1624 => x"53776170",
  1625 => x"206a6f79",
  1626 => x"3a204f6e",
  1627 => x"00000000",
  1628 => x"5363616e",
  1629 => x"6c696e65",
  1630 => x"733a204e",
  1631 => x"6f6e6500",
  1632 => x"5363616e",
  1633 => x"4c696e65",
  1634 => x"733a2048",
  1635 => x"51327800",
  1636 => x"5363616e",
  1637 => x"6c696e65",
  1638 => x"733a2043",
  1639 => x"52542032",
  1640 => x"35250000",
  1641 => x"5363616e",
  1642 => x"6c696e65",
  1643 => x"733a2043",
  1644 => x"52542035",
  1645 => x"30250000",
  1646 => x"5363616e",
  1647 => x"6c696e65",
  1648 => x"733a2043",
  1649 => x"52542037",
  1650 => x"35250000",
  1651 => x"43617267",
  1652 => x"61204661",
  1653 => x"6c6c6964",
  1654 => x"61000000",
  1655 => x"4f4b0000",
  1656 => x"16200000",
  1657 => x"14200000",
  1658 => x"15200000",
  1659 => x"53442069",
  1660 => x"6e69742e",
  1661 => x"2e2e0a00",
  1662 => x"53442063",
  1663 => x"61726420",
  1664 => x"72657365",
  1665 => x"74206661",
  1666 => x"696c6564",
  1667 => x"210a0000",
  1668 => x"53444843",
  1669 => x"20657272",
  1670 => x"6f72210a",
  1671 => x"00000000",
  1672 => x"57726974",
  1673 => x"65206661",
  1674 => x"696c6564",
  1675 => x"0a000000",
  1676 => x"52656164",
  1677 => x"20666169",
  1678 => x"6c65640a",
  1679 => x"00000000",
  1680 => x"43617264",
  1681 => x"20696e69",
  1682 => x"74206661",
  1683 => x"696c6564",
  1684 => x"0a000000",
  1685 => x"46415431",
  1686 => x"36202020",
  1687 => x"00000000",
  1688 => x"46415433",
  1689 => x"32202020",
  1690 => x"00000000",
  1691 => x"4e6f2070",
  1692 => x"61727469",
  1693 => x"74696f6e",
  1694 => x"20736967",
  1695 => x"0a000000",
  1696 => x"42616420",
  1697 => x"70617274",
  1698 => x"0a000000",
  1699 => x"4261636b",
  1700 => x"00000000",
  1701 => x"00000002",
  1702 => x"00000002",
  1703 => x"000017f8",
  1704 => x"00000000",
  1705 => x"00000002",
  1706 => x"00001810",
  1707 => x"00000000",
  1708 => x"00000002",
  1709 => x"00001828",
  1710 => x"0000034e",
  1711 => x"00000003",
  1712 => x"00001b54",
  1713 => x"00000004",
  1714 => x"00000003",
  1715 => x"00001b4c",
  1716 => x"00000002",
  1717 => x"00000003",
  1718 => x"00001b44",
  1719 => x"00000002",
  1720 => x"00000003",
  1721 => x"00001b24",
  1722 => x"00000008",
  1723 => x"00000003",
  1724 => x"00001b1c",
  1725 => x"00000002",
  1726 => x"00000002",
  1727 => x"00001830",
  1728 => x"000017c2",
  1729 => x"00000002",
  1730 => x"00001848",
  1731 => x"000006c1",
  1732 => x"00000000",
  1733 => x"00000000",
  1734 => x"00000000",
  1735 => x"00001850",
  1736 => x"00001864",
  1737 => x"00001878",
  1738 => x"00001888",
  1739 => x"000018a0",
  1740 => x"000018b8",
  1741 => x"000018d0",
  1742 => x"000018e8",
  1743 => x"00001900",
  1744 => x"00001918",
  1745 => x"00001930",
  1746 => x"00001940",
  1747 => x"00001950",
  1748 => x"00001960",
  1749 => x"00001970",
  1750 => x"00001980",
  1751 => x"00001990",
  1752 => x"000019a4",
  1753 => x"000019b8",
  1754 => x"00000004",
  1755 => x"000019cc",
  1756 => x"00001b68",
  1757 => x"00000004",
  1758 => x"000019dc",
  1759 => x"00001a98",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000000",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"00000000",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"00000002",
  1785 => x"00002040",
  1786 => x"000015bb",
  1787 => x"00000002",
  1788 => x"0000205e",
  1789 => x"000015bb",
  1790 => x"00000002",
  1791 => x"0000207c",
  1792 => x"000015bb",
  1793 => x"00000002",
  1794 => x"0000209a",
  1795 => x"000015bb",
  1796 => x"00000002",
  1797 => x"000020b8",
  1798 => x"000015bb",
  1799 => x"00000002",
  1800 => x"000020d6",
  1801 => x"000015bb",
  1802 => x"00000002",
  1803 => x"000020f4",
  1804 => x"000015bb",
  1805 => x"00000002",
  1806 => x"00002112",
  1807 => x"000015bb",
  1808 => x"00000002",
  1809 => x"00002130",
  1810 => x"000015bb",
  1811 => x"00000002",
  1812 => x"0000214e",
  1813 => x"000015bb",
  1814 => x"00000002",
  1815 => x"0000216c",
  1816 => x"000015bb",
  1817 => x"00000002",
  1818 => x"0000218a",
  1819 => x"000015bb",
  1820 => x"00000002",
  1821 => x"000021a8",
  1822 => x"000015bb",
  1823 => x"00000004",
  1824 => x"00001a8c",
  1825 => x"00000000",
  1826 => x"00000000",
  1827 => x"00000000",
  1828 => x"00001756",
  1829 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

