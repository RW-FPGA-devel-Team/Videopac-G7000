-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d1",
     9 => x"9c080b0b",
    10 => x"80d1a008",
    11 => x"0b0b80d1",
    12 => x"a4080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d1a40c0b",
    16 => x"0b80d1a0",
    17 => x"0c0b0b80",
    18 => x"d19c0c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbd98",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d19c70",
    57 => x"80dbd827",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518aa2",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d1",
    65 => x"ac0c9f0b",
    66 => x"80d1b00c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d1b008ff",
    70 => x"0580d1b0",
    71 => x"0c80d1b0",
    72 => x"088025e8",
    73 => x"3880d1ac",
    74 => x"08ff0580",
    75 => x"d1ac0c80",
    76 => x"d1ac0880",
    77 => x"25d03880",
    78 => x"0b80d1b0",
    79 => x"0c800b80",
    80 => x"d1ac0c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d1ac08",
   100 => x"25913882",
   101 => x"c82d80d1",
   102 => x"ac08ff05",
   103 => x"80d1ac0c",
   104 => x"838a0480",
   105 => x"d1ac0880",
   106 => x"d1b00853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d1ac08",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d1b00881",
   116 => x"0580d1b0",
   117 => x"0c80d1b0",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d1b0",
   121 => x"0c80d1ac",
   122 => x"08810580",
   123 => x"d1ac0c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d1",
   128 => x"b0088105",
   129 => x"80d1b00c",
   130 => x"80d1b008",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d1b0",
   134 => x"0c80d1ac",
   135 => x"08810580",
   136 => x"d1ac0c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d1b40cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d1b40c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d1",
   177 => x"b4088407",
   178 => x"80d1b40c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5485bc74",
   182 => x"258f3882",
   183 => x"0b0b0b80",
   184 => x"c8d40c80",
   185 => x"d05385f3",
   186 => x"04810b0b",
   187 => x"0b80c8d4",
   188 => x"0cbc530b",
   189 => x"0b80c8d4",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0cfc0875",
   193 => x"7531ffb0",
   194 => x"05ff1371",
   195 => x"712cff94",
   196 => x"1a709f2a",
   197 => x"1170812c",
   198 => x"80d1b408",
   199 => x"52545153",
   200 => x"57535152",
   201 => x"5276802e",
   202 => x"85387081",
   203 => x"075170f6",
   204 => x"940c7209",
   205 => x"8105f680",
   206 => x"0c710981",
   207 => x"05f6840c",
   208 => x"0294050d",
   209 => x"0402f405",
   210 => x"0d745372",
   211 => x"70810554",
   212 => x"80f52d52",
   213 => x"71802e89",
   214 => x"38715183",
   215 => x"842d86cb",
   216 => x"04810b80",
   217 => x"d19c0c02",
   218 => x"8c050d04",
   219 => x"02fc050d",
   220 => x"81808051",
   221 => x"c0115170",
   222 => x"fb380284",
   223 => x"050d0402",
   224 => x"fc050dec",
   225 => x"5183710c",
   226 => x"86ec2d82",
   227 => x"710c0284",
   228 => x"050d0402",
   229 => x"fc050d84",
   230 => x"bf5186ec",
   231 => x"2dff1151",
   232 => x"708025f6",
   233 => x"38028405",
   234 => x"0d040402",
   235 => x"fc050d92",
   236 => x"a62d80d1",
   237 => x"9c0880ce",
   238 => x"d80c80cd",
   239 => x"b45194de",
   240 => x"2d028405",
   241 => x"0d0402fc",
   242 => x"050d92a6",
   243 => x"2d80d19c",
   244 => x"0880cda4",
   245 => x"0c80cc80",
   246 => x"5194de2d",
   247 => x"0284050d",
   248 => x"0402dc05",
   249 => x"0d7a5580",
   250 => x"59840bec",
   251 => x"0c80c8dc",
   252 => x"085380c8",
   253 => x"d808812e",
   254 => x"0981068c",
   255 => x"38728280",
   256 => x"0780c8dc",
   257 => x"0c889304",
   258 => x"72828007",
   259 => x"82803280",
   260 => x"c8dc0c80",
   261 => x"c8dc08fc",
   262 => x"0c86ec2d",
   263 => x"745280d1",
   264 => x"b851b3d5",
   265 => x"2d80d19c",
   266 => x"08802e81",
   267 => x"ae3880d1",
   268 => x"bc085480",
   269 => x"5673852e",
   270 => x"098106a5",
   271 => x"38745186",
   272 => x"c52d8793",
   273 => x"2d87932d",
   274 => x"87932d87",
   275 => x"932d8793",
   276 => x"2d87932d",
   277 => x"80d1c408",
   278 => x"5194de2d",
   279 => x"81538a98",
   280 => x"0473f80c",
   281 => x"a50bec0c",
   282 => x"87932d84",
   283 => x"0bec0c75",
   284 => x"ff155758",
   285 => x"75802e8b",
   286 => x"38811876",
   287 => x"812a5758",
   288 => x"88f404f7",
   289 => x"18588159",
   290 => x"80742580",
   291 => x"ce387752",
   292 => x"755184a8",
   293 => x"2d80d290",
   294 => x"5280d1b8",
   295 => x"51b6a22d",
   296 => x"80d19c08",
   297 => x"802e9b38",
   298 => x"80d29057",
   299 => x"83fc5576",
   300 => x"70840558",
   301 => x"08e80cfc",
   302 => x"15557480",
   303 => x"25f13889",
   304 => x"ca0480d1",
   305 => x"9c085984",
   306 => x"805480d1",
   307 => x"b851b5f2",
   308 => x"2dfc8014",
   309 => x"81175754",
   310 => x"89880480",
   311 => x"c8d80853",
   312 => x"72893872",
   313 => x"5186ff2d",
   314 => x"8a820480",
   315 => x"0b80c8d8",
   316 => x"0c80c8dc",
   317 => x"08828007",
   318 => x"82803270",
   319 => x"80c8dc0c",
   320 => x"fc0c7880",
   321 => x"2e893880",
   322 => x"d1c40851",
   323 => x"8a930480",
   324 => x"cbdc5194",
   325 => x"de2d7853",
   326 => x"7280d19c",
   327 => x"0c02a405",
   328 => x"0d0402ec",
   329 => x"050d900b",
   330 => x"80c8dc0c",
   331 => x"805186ff",
   332 => x"2d840bec",
   333 => x"0c91f62d",
   334 => x"8ea12d81",
   335 => x"f92d8353",
   336 => x"91d92d81",
   337 => x"51858d2d",
   338 => x"ff135372",
   339 => x"8025f138",
   340 => x"840bec0c",
   341 => x"80c78851",
   342 => x"86c52daa",
   343 => x"8d2d80d1",
   344 => x"9c08802e",
   345 => x"83a43881",
   346 => x"0bec0c84",
   347 => x"0bec0cbd",
   348 => x"a85280d1",
   349 => x"b851b3d5",
   350 => x"2d80d19c",
   351 => x"08802e80",
   352 => x"cb3880d2",
   353 => x"905280d1",
   354 => x"b851b6a2",
   355 => x"2d80d19c",
   356 => x"08802eb8",
   357 => x"3880d290",
   358 => x"0b80f52d",
   359 => x"80cfc80c",
   360 => x"80d2910b",
   361 => x"80f52d80",
   362 => x"cfcc0c80",
   363 => x"d2920b80",
   364 => x"f52d80cf",
   365 => x"d00c80d2",
   366 => x"930b80f5",
   367 => x"2d80cfd4",
   368 => x"0c80d294",
   369 => x"0b80f52d",
   370 => x"80cfd80c",
   371 => x"bdb85280",
   372 => x"d1b851b3",
   373 => x"d52d80d1",
   374 => x"9c08802e",
   375 => x"80cb3880",
   376 => x"d2905280",
   377 => x"d1b851b6",
   378 => x"a22d80d1",
   379 => x"9c08802e",
   380 => x"b83880d2",
   381 => x"900b80f5",
   382 => x"2d80cfb4",
   383 => x"0c80d291",
   384 => x"0b80f52d",
   385 => x"80cfb80c",
   386 => x"80d2920b",
   387 => x"80f52d80",
   388 => x"cfbc0c80",
   389 => x"d2930b80",
   390 => x"f52d80cf",
   391 => x"c00c80d2",
   392 => x"940b80f5",
   393 => x"2d80cfc4",
   394 => x"0c87e151",
   395 => x"bd922d80",
   396 => x"c8dc0880",
   397 => x"cfb00c80",
   398 => x"c8dc08fc",
   399 => x"0c80d1f0",
   400 => x"08882a70",
   401 => x"81065153",
   402 => x"72802e8c",
   403 => x"3880caa8",
   404 => x"0b80d1c4",
   405 => x"0c8ce004",
   406 => x"80c8e00b",
   407 => x"80d1c40c",
   408 => x"80d1c408",
   409 => x"5194de2d",
   410 => x"860b80d2",
   411 => x"840c92af",
   412 => x"2d8ead2d",
   413 => x"94f12d80",
   414 => x"d1c40880",
   415 => x"e81180f5",
   416 => x"2d70842b",
   417 => x"7080c8dc",
   418 => x"0c80f413",
   419 => x"80f52d70",
   420 => x"852b7207",
   421 => x"7080c8dc",
   422 => x"0c818015",
   423 => x"80f52d70",
   424 => x"892b7207",
   425 => x"7080c8dc",
   426 => x"0c80cfb0",
   427 => x"08708106",
   428 => x"53535355",
   429 => x"52525656",
   430 => x"5372802e",
   431 => x"88387481",
   432 => x"0780c8dc",
   433 => x"0c73812a",
   434 => x"70810651",
   435 => x"5372802e",
   436 => x"8b3880c8",
   437 => x"dc088207",
   438 => x"80c8dc0c",
   439 => x"73822a70",
   440 => x"81065153",
   441 => x"72802e8c",
   442 => x"3880c8dc",
   443 => x"08818007",
   444 => x"80c8dc0c",
   445 => x"80c8dc08",
   446 => x"fc0c8653",
   447 => x"80d19c08",
   448 => x"83388453",
   449 => x"72ec0c8c",
   450 => x"f104800b",
   451 => x"80d19c0c",
   452 => x"0294050d",
   453 => x"0471980c",
   454 => x"04ffb008",
   455 => x"80d19c0c",
   456 => x"04810bff",
   457 => x"b00c0480",
   458 => x"0bffb00c",
   459 => x"0402f405",
   460 => x"0d8fbb04",
   461 => x"80d19c08",
   462 => x"81f02e09",
   463 => x"81068a38",
   464 => x"810b80cf",
   465 => x"a80c8fbb",
   466 => x"0480d19c",
   467 => x"0881e02e",
   468 => x"0981068a",
   469 => x"38810b80",
   470 => x"cfac0c8f",
   471 => x"bb0480d1",
   472 => x"9c085280",
   473 => x"cfac0880",
   474 => x"2e893880",
   475 => x"d19c0881",
   476 => x"80055271",
   477 => x"842c728f",
   478 => x"06535380",
   479 => x"cfa80880",
   480 => x"2e9a3872",
   481 => x"842980ce",
   482 => x"e8057213",
   483 => x"81712b70",
   484 => x"09730806",
   485 => x"730c5153",
   486 => x"538faf04",
   487 => x"72842980",
   488 => x"cee80572",
   489 => x"1383712b",
   490 => x"72080772",
   491 => x"0c535380",
   492 => x"0b80cfac",
   493 => x"0c800b80",
   494 => x"cfa80c80",
   495 => x"d1c85190",
   496 => x"c22d80d1",
   497 => x"9c08ff24",
   498 => x"feea3880",
   499 => x"0b80d19c",
   500 => x"0c028c05",
   501 => x"0d0402f8",
   502 => x"050d80ce",
   503 => x"e8528f51",
   504 => x"80727084",
   505 => x"05540cff",
   506 => x"11517080",
   507 => x"25f23802",
   508 => x"88050d04",
   509 => x"02f0050d",
   510 => x"75518ea7",
   511 => x"2d70822c",
   512 => x"fc0680ce",
   513 => x"e8117210",
   514 => x"9e067108",
   515 => x"70722a70",
   516 => x"83068274",
   517 => x"2b700974",
   518 => x"06760c54",
   519 => x"51565753",
   520 => x"51538ea1",
   521 => x"2d7180d1",
   522 => x"9c0c0290",
   523 => x"050d0402",
   524 => x"fc050d72",
   525 => x"5180710c",
   526 => x"800b8412",
   527 => x"0c028405",
   528 => x"0d0402f0",
   529 => x"050d7570",
   530 => x"08841208",
   531 => x"535353ff",
   532 => x"5471712e",
   533 => x"a8388ea7",
   534 => x"2d841308",
   535 => x"70842914",
   536 => x"88117008",
   537 => x"7081ff06",
   538 => x"84180881",
   539 => x"11870684",
   540 => x"1a0c5351",
   541 => x"55515151",
   542 => x"8ea12d71",
   543 => x"547380d1",
   544 => x"9c0c0290",
   545 => x"050d0402",
   546 => x"f4050d8e",
   547 => x"a72de008",
   548 => x"708b2a70",
   549 => x"81065152",
   550 => x"5370802e",
   551 => x"a13880d1",
   552 => x"c8087084",
   553 => x"2980d1d0",
   554 => x"057481ff",
   555 => x"06710c51",
   556 => x"5180d1c8",
   557 => x"08811187",
   558 => x"0680d1c8",
   559 => x"0c51728c",
   560 => x"2c83ff06",
   561 => x"80d1f00c",
   562 => x"800b80d1",
   563 => x"f40c8e99",
   564 => x"2d8ea12d",
   565 => x"028c050d",
   566 => x"0402fc05",
   567 => x"0d8ea72d",
   568 => x"810b80d1",
   569 => x"f40c8ea1",
   570 => x"2d80d1f4",
   571 => x"085170f9",
   572 => x"38028405",
   573 => x"0d0402fc",
   574 => x"050d80d1",
   575 => x"c85190af",
   576 => x"2d8fd62d",
   577 => x"9187518e",
   578 => x"952d0284",
   579 => x"050d0402",
   580 => x"fc050d8f",
   581 => x"cf5186ec",
   582 => x"2dff1151",
   583 => x"708025f6",
   584 => x"38028405",
   585 => x"0d0480d1",
   586 => x"fc0880d1",
   587 => x"9c0c0402",
   588 => x"fc050d81",
   589 => x"0b80cfdc",
   590 => x"0c815185",
   591 => x"8d2d0284",
   592 => x"050d0402",
   593 => x"fc050d92",
   594 => x"cd048ead",
   595 => x"2d80f651",
   596 => x"8ff42d80",
   597 => x"d19c08f2",
   598 => x"3880da51",
   599 => x"8ff42d80",
   600 => x"d19c08e6",
   601 => x"3880cfd8",
   602 => x"08518ff4",
   603 => x"2d80d19c",
   604 => x"08d83880",
   605 => x"d19c0880",
   606 => x"cfdc0c80",
   607 => x"d19c0851",
   608 => x"858d2d02",
   609 => x"84050d04",
   610 => x"02ec050d",
   611 => x"76548052",
   612 => x"870b8815",
   613 => x"80f52d56",
   614 => x"53747224",
   615 => x"8338a053",
   616 => x"72518384",
   617 => x"2d81128b",
   618 => x"1580f52d",
   619 => x"54527272",
   620 => x"25de3802",
   621 => x"94050d04",
   622 => x"02f0050d",
   623 => x"80d1fc08",
   624 => x"5481f92d",
   625 => x"800b80d2",
   626 => x"800c7308",
   627 => x"802e8189",
   628 => x"38820b80",
   629 => x"d1b00c80",
   630 => x"d280088f",
   631 => x"0680d1ac",
   632 => x"0c730852",
   633 => x"71832e96",
   634 => x"38718326",
   635 => x"89387181",
   636 => x"2eb03894",
   637 => x"c2047185",
   638 => x"2ea03894",
   639 => x"c2048814",
   640 => x"80f52d84",
   641 => x"150880c7",
   642 => x"a0535452",
   643 => x"86c52d71",
   644 => x"84291370",
   645 => x"08525294",
   646 => x"c6047351",
   647 => x"93882d94",
   648 => x"c20480cf",
   649 => x"b0088815",
   650 => x"082c7081",
   651 => x"06515271",
   652 => x"802e8838",
   653 => x"80c7a451",
   654 => x"94bf0480",
   655 => x"c7a85186",
   656 => x"c52d8414",
   657 => x"085186c5",
   658 => x"2d80d280",
   659 => x"08810580",
   660 => x"d2800c8c",
   661 => x"145493ca",
   662 => x"04029005",
   663 => x"0d047180",
   664 => x"d1fc0c93",
   665 => x"b82d80d2",
   666 => x"8008ff05",
   667 => x"80d2840c",
   668 => x"0402e805",
   669 => x"0d80d1fc",
   670 => x"0880d288",
   671 => x"08575580",
   672 => x"f6518ff4",
   673 => x"2d80d19c",
   674 => x"08812a70",
   675 => x"81065152",
   676 => x"71802ea2",
   677 => x"38959b04",
   678 => x"8ead2d80",
   679 => x"f6518ff4",
   680 => x"2d80d19c",
   681 => x"08f23880",
   682 => x"cfdc0881",
   683 => x"327080cf",
   684 => x"dc0c5185",
   685 => x"8d2d800b",
   686 => x"80d1f80c",
   687 => x"86518ff4",
   688 => x"2d80d19c",
   689 => x"08812a70",
   690 => x"81065152",
   691 => x"71802e8b",
   692 => x"3880c8dc",
   693 => x"08903280",
   694 => x"c8dc0c8c",
   695 => x"518ff42d",
   696 => x"80d19c08",
   697 => x"812a7081",
   698 => x"06515271",
   699 => x"802e80d1",
   700 => x"3880cfb4",
   701 => x"0880cfc8",
   702 => x"0880cfb4",
   703 => x"0c80cfc8",
   704 => x"0c80cfb8",
   705 => x"0880cfcc",
   706 => x"0880cfb8",
   707 => x"0c80cfcc",
   708 => x"0c80cfbc",
   709 => x"0880cfd0",
   710 => x"0880cfbc",
   711 => x"0c80cfd0",
   712 => x"0c80cfc0",
   713 => x"0880cfd4",
   714 => x"0880cfc0",
   715 => x"0c80cfd4",
   716 => x"0c80cfc4",
   717 => x"0880cfd8",
   718 => x"0880cfc4",
   719 => x"0c80cfd8",
   720 => x"0c80d1f0",
   721 => x"08a00652",
   722 => x"80722596",
   723 => x"38928f2d",
   724 => x"8ead2d80",
   725 => x"cfdc0881",
   726 => x"327080cf",
   727 => x"dc0c5185",
   728 => x"8d2d80cf",
   729 => x"dc0882ef",
   730 => x"3880cfc8",
   731 => x"08518ff4",
   732 => x"2d80d19c",
   733 => x"08802e8b",
   734 => x"3880d1f8",
   735 => x"08810780",
   736 => x"d1f80c80",
   737 => x"cfcc0851",
   738 => x"8ff42d80",
   739 => x"d19c0880",
   740 => x"2e8b3880",
   741 => x"d1f80882",
   742 => x"0780d1f8",
   743 => x"0c80cfd0",
   744 => x"08518ff4",
   745 => x"2d80d19c",
   746 => x"08802e8b",
   747 => x"3880d1f8",
   748 => x"08840780",
   749 => x"d1f80c80",
   750 => x"cfd40851",
   751 => x"8ff42d80",
   752 => x"d19c0880",
   753 => x"2e8b3880",
   754 => x"d1f80888",
   755 => x"0780d1f8",
   756 => x"0c80cfd8",
   757 => x"08518ff4",
   758 => x"2d80d19c",
   759 => x"08802e8b",
   760 => x"3880d1f8",
   761 => x"08900780",
   762 => x"d1f80c80",
   763 => x"cfb40851",
   764 => x"8ff42d80",
   765 => x"d19c0880",
   766 => x"2e8c3880",
   767 => x"d1f80882",
   768 => x"800780d1",
   769 => x"f80c80cf",
   770 => x"b808518f",
   771 => x"f42d80d1",
   772 => x"9c08802e",
   773 => x"8c3880d1",
   774 => x"f8088480",
   775 => x"0780d1f8",
   776 => x"0c80cfbc",
   777 => x"08518ff4",
   778 => x"2d80d19c",
   779 => x"08802e8c",
   780 => x"3880d1f8",
   781 => x"08888007",
   782 => x"80d1f80c",
   783 => x"80cfc008",
   784 => x"518ff42d",
   785 => x"80d19c08",
   786 => x"802e8c38",
   787 => x"80d1f808",
   788 => x"90800780",
   789 => x"d1f80c80",
   790 => x"cfc40851",
   791 => x"8ff42d80",
   792 => x"d19c0880",
   793 => x"2e8c3880",
   794 => x"d1f808a0",
   795 => x"800780d1",
   796 => x"f80c9451",
   797 => x"8ff42d80",
   798 => x"d19c0852",
   799 => x"91518ff4",
   800 => x"2d7180d1",
   801 => x"9c080652",
   802 => x"80e6518f",
   803 => x"f42d7180",
   804 => x"d19c0806",
   805 => x"5271802e",
   806 => x"8d3880d1",
   807 => x"f8088480",
   808 => x"800780d1",
   809 => x"f80c80fe",
   810 => x"518ff42d",
   811 => x"80d19c08",
   812 => x"5287518f",
   813 => x"f42d7180",
   814 => x"d19c0807",
   815 => x"5271802e",
   816 => x"8d3880d1",
   817 => x"f8088880",
   818 => x"800780d1",
   819 => x"f80c80d1",
   820 => x"f808ed0c",
   821 => x"a1e20494",
   822 => x"518ff42d",
   823 => x"80d19c08",
   824 => x"5291518f",
   825 => x"f42d7180",
   826 => x"d19c0806",
   827 => x"5280e651",
   828 => x"8ff42d71",
   829 => x"80d19c08",
   830 => x"06527180",
   831 => x"2e8d3880",
   832 => x"d1f80884",
   833 => x"80800780",
   834 => x"d1f80c80",
   835 => x"fe518ff4",
   836 => x"2d80d19c",
   837 => x"08528751",
   838 => x"8ff42d71",
   839 => x"80d19c08",
   840 => x"07527180",
   841 => x"2e8d3880",
   842 => x"d1f80888",
   843 => x"80800780",
   844 => x"d1f80c80",
   845 => x"d1f808ed",
   846 => x"0c81f551",
   847 => x"8ff42d80",
   848 => x"d19c0881",
   849 => x"2a708106",
   850 => x"515271a4",
   851 => x"3880cfc8",
   852 => x"08518ff4",
   853 => x"2d80d19c",
   854 => x"08812a70",
   855 => x"81065152",
   856 => x"718e3880",
   857 => x"d1f00881",
   858 => x"06528072",
   859 => x"2580c238",
   860 => x"80d1f008",
   861 => x"81065280",
   862 => x"72258438",
   863 => x"928f2d80",
   864 => x"d2840852",
   865 => x"71802e8a",
   866 => x"38ff1280",
   867 => x"d2840c9b",
   868 => x"b10480d2",
   869 => x"80081080",
   870 => x"d2800805",
   871 => x"70842916",
   872 => x"51528812",
   873 => x"08802e89",
   874 => x"38ff5188",
   875 => x"12085271",
   876 => x"2d81f251",
   877 => x"8ff42d80",
   878 => x"d19c0881",
   879 => x"2a708106",
   880 => x"515271a4",
   881 => x"3880cfcc",
   882 => x"08518ff4",
   883 => x"2d80d19c",
   884 => x"08812a70",
   885 => x"81065152",
   886 => x"718e3880",
   887 => x"d1f00882",
   888 => x"06528072",
   889 => x"2580c338",
   890 => x"80d1f008",
   891 => x"82065280",
   892 => x"72258438",
   893 => x"928f2d80",
   894 => x"d28008ff",
   895 => x"1180d284",
   896 => x"08565353",
   897 => x"7372258a",
   898 => x"38811480",
   899 => x"d2840c9c",
   900 => x"aa047210",
   901 => x"13708429",
   902 => x"16515288",
   903 => x"1208802e",
   904 => x"8938fe51",
   905 => x"88120852",
   906 => x"712d81fd",
   907 => x"518ff42d",
   908 => x"80d19c08",
   909 => x"812a7081",
   910 => x"06515271",
   911 => x"a43880cf",
   912 => x"d008518f",
   913 => x"f42d80d1",
   914 => x"9c08812a",
   915 => x"70810651",
   916 => x"52718e38",
   917 => x"80d1f008",
   918 => x"84065280",
   919 => x"722580c0",
   920 => x"3880d1f0",
   921 => x"08840652",
   922 => x"80722584",
   923 => x"38928f2d",
   924 => x"80d28408",
   925 => x"802e8a38",
   926 => x"800b80d2",
   927 => x"840c9da0",
   928 => x"0480d280",
   929 => x"081080d2",
   930 => x"80080570",
   931 => x"84291651",
   932 => x"52881208",
   933 => x"802e8938",
   934 => x"fd518812",
   935 => x"0852712d",
   936 => x"81fa518f",
   937 => x"f42d80d1",
   938 => x"9c08812a",
   939 => x"70810651",
   940 => x"5271a438",
   941 => x"80cfd408",
   942 => x"518ff42d",
   943 => x"80d19c08",
   944 => x"812a7081",
   945 => x"06515271",
   946 => x"8e3880d1",
   947 => x"f0088806",
   948 => x"52807225",
   949 => x"80c03880",
   950 => x"d1f00888",
   951 => x"06528072",
   952 => x"25843892",
   953 => x"8f2d80d2",
   954 => x"8008ff11",
   955 => x"545280d2",
   956 => x"84087325",
   957 => x"89387280",
   958 => x"d2840c9e",
   959 => x"96047110",
   960 => x"12708429",
   961 => x"16515288",
   962 => x"1208802e",
   963 => x"8938fc51",
   964 => x"88120852",
   965 => x"712d80d2",
   966 => x"84087053",
   967 => x"5473802e",
   968 => x"8a388c15",
   969 => x"ff155555",
   970 => x"9e9d0482",
   971 => x"0b80d1b0",
   972 => x"0c718f06",
   973 => x"80d1ac0c",
   974 => x"81eb518f",
   975 => x"f42d80d1",
   976 => x"9c08812a",
   977 => x"70810651",
   978 => x"5271802e",
   979 => x"ad387408",
   980 => x"852e0981",
   981 => x"06a43888",
   982 => x"1580f52d",
   983 => x"ff055271",
   984 => x"881681b7",
   985 => x"2d71982b",
   986 => x"52718025",
   987 => x"8838800b",
   988 => x"881681b7",
   989 => x"2d745193",
   990 => x"882d81f4",
   991 => x"518ff42d",
   992 => x"80d19c08",
   993 => x"812a7081",
   994 => x"06515271",
   995 => x"802eb338",
   996 => x"7408852e",
   997 => x"098106aa",
   998 => x"38881580",
   999 => x"f52d8105",
  1000 => x"52718816",
  1001 => x"81b72d71",
  1002 => x"81ff068b",
  1003 => x"1680f52d",
  1004 => x"54527272",
  1005 => x"27873872",
  1006 => x"881681b7",
  1007 => x"2d745193",
  1008 => x"882d80da",
  1009 => x"518ff42d",
  1010 => x"80d19c08",
  1011 => x"812a7081",
  1012 => x"06515271",
  1013 => x"8e3880d1",
  1014 => x"f0089006",
  1015 => x"52807225",
  1016 => x"81bc3880",
  1017 => x"d1fc0880",
  1018 => x"d1f00890",
  1019 => x"06535380",
  1020 => x"72258438",
  1021 => x"928f2d80",
  1022 => x"d2840854",
  1023 => x"73802e8a",
  1024 => x"388c13ff",
  1025 => x"1555539f",
  1026 => x"fc047208",
  1027 => x"5271822e",
  1028 => x"a6387182",
  1029 => x"26893871",
  1030 => x"812eaa38",
  1031 => x"a19e0471",
  1032 => x"832eb438",
  1033 => x"71842e09",
  1034 => x"810680f2",
  1035 => x"38881308",
  1036 => x"5194de2d",
  1037 => x"a19e0480",
  1038 => x"d2840851",
  1039 => x"88130852",
  1040 => x"712da19e",
  1041 => x"04810b88",
  1042 => x"14082b80",
  1043 => x"cfb00832",
  1044 => x"80cfb00c",
  1045 => x"a0f20488",
  1046 => x"1380f52d",
  1047 => x"81058b14",
  1048 => x"80f52d53",
  1049 => x"54717424",
  1050 => x"83388054",
  1051 => x"73881481",
  1052 => x"b72d93b8",
  1053 => x"2da19e04",
  1054 => x"7508802e",
  1055 => x"a4387508",
  1056 => x"518ff42d",
  1057 => x"80d19c08",
  1058 => x"81065271",
  1059 => x"802e8c38",
  1060 => x"80d28408",
  1061 => x"51841608",
  1062 => x"52712d88",
  1063 => x"165675d8",
  1064 => x"38805480",
  1065 => x"0b80d1b0",
  1066 => x"0c738f06",
  1067 => x"80d1ac0c",
  1068 => x"a0527380",
  1069 => x"d284082e",
  1070 => x"09810699",
  1071 => x"3880d280",
  1072 => x"08ff0574",
  1073 => x"32700981",
  1074 => x"05707207",
  1075 => x"9f2a9171",
  1076 => x"31515153",
  1077 => x"53715183",
  1078 => x"842d8114",
  1079 => x"548e7425",
  1080 => x"c23880cf",
  1081 => x"dc0880d1",
  1082 => x"9c0c0298",
  1083 => x"050d0402",
  1084 => x"f4050dd4",
  1085 => x"5281ff72",
  1086 => x"0c710853",
  1087 => x"81ff720c",
  1088 => x"72882b83",
  1089 => x"fe800672",
  1090 => x"087081ff",
  1091 => x"06515253",
  1092 => x"81ff720c",
  1093 => x"72710788",
  1094 => x"2b720870",
  1095 => x"81ff0651",
  1096 => x"525381ff",
  1097 => x"720c7271",
  1098 => x"07882b72",
  1099 => x"087081ff",
  1100 => x"06720780",
  1101 => x"d19c0c52",
  1102 => x"53028c05",
  1103 => x"0d0402f4",
  1104 => x"050d7476",
  1105 => x"7181ff06",
  1106 => x"d40c5353",
  1107 => x"80d28c08",
  1108 => x"85387189",
  1109 => x"2b527198",
  1110 => x"2ad40c71",
  1111 => x"902a7081",
  1112 => x"ff06d40c",
  1113 => x"5171882a",
  1114 => x"7081ff06",
  1115 => x"d40c5171",
  1116 => x"81ff06d4",
  1117 => x"0c72902a",
  1118 => x"7081ff06",
  1119 => x"d40c51d4",
  1120 => x"087081ff",
  1121 => x"06515182",
  1122 => x"b8bf5270",
  1123 => x"81ff2e09",
  1124 => x"81069438",
  1125 => x"81ff0bd4",
  1126 => x"0cd40870",
  1127 => x"81ff06ff",
  1128 => x"14545151",
  1129 => x"71e53870",
  1130 => x"80d19c0c",
  1131 => x"028c050d",
  1132 => x"0402fc05",
  1133 => x"0d81c751",
  1134 => x"81ff0bd4",
  1135 => x"0cff1151",
  1136 => x"708025f4",
  1137 => x"38028405",
  1138 => x"0d0402f4",
  1139 => x"050d81ff",
  1140 => x"0bd40c93",
  1141 => x"53805287",
  1142 => x"fc80c151",
  1143 => x"a2be2d80",
  1144 => x"d19c088b",
  1145 => x"3881ff0b",
  1146 => x"d40c8153",
  1147 => x"a3f804a3",
  1148 => x"b12dff13",
  1149 => x"5372de38",
  1150 => x"7280d19c",
  1151 => x"0c028c05",
  1152 => x"0d0402ec",
  1153 => x"050d810b",
  1154 => x"80d28c0c",
  1155 => x"8454d008",
  1156 => x"708f2a70",
  1157 => x"81065151",
  1158 => x"5372f338",
  1159 => x"72d00ca3",
  1160 => x"b12d80c7",
  1161 => x"ac5186c5",
  1162 => x"2dd00870",
  1163 => x"8f2a7081",
  1164 => x"06515153",
  1165 => x"72f33881",
  1166 => x"0bd00cb1",
  1167 => x"53805284",
  1168 => x"d480c051",
  1169 => x"a2be2d80",
  1170 => x"d19c0881",
  1171 => x"2e933872",
  1172 => x"822ebf38",
  1173 => x"ff135372",
  1174 => x"e438ff14",
  1175 => x"5473ffae",
  1176 => x"38a3b12d",
  1177 => x"83aa5284",
  1178 => x"9c80c851",
  1179 => x"a2be2d80",
  1180 => x"d19c0881",
  1181 => x"2e098106",
  1182 => x"9338a1ef",
  1183 => x"2d80d19c",
  1184 => x"0883ffff",
  1185 => x"06537283",
  1186 => x"aa2e9f38",
  1187 => x"a3ca2da5",
  1188 => x"a50480c7",
  1189 => x"b85186c5",
  1190 => x"2d8053a6",
  1191 => x"fa0480c7",
  1192 => x"d05186c5",
  1193 => x"2d8054a6",
  1194 => x"cb0481ff",
  1195 => x"0bd40cb1",
  1196 => x"54a3b12d",
  1197 => x"8fcf5380",
  1198 => x"5287fc80",
  1199 => x"f751a2be",
  1200 => x"2d80d19c",
  1201 => x"085580d1",
  1202 => x"9c08812e",
  1203 => x"0981069c",
  1204 => x"3881ff0b",
  1205 => x"d40c820a",
  1206 => x"52849c80",
  1207 => x"e951a2be",
  1208 => x"2d80d19c",
  1209 => x"08802e8d",
  1210 => x"38a3b12d",
  1211 => x"ff135372",
  1212 => x"c638a6be",
  1213 => x"0481ff0b",
  1214 => x"d40c80d1",
  1215 => x"9c085287",
  1216 => x"fc80fa51",
  1217 => x"a2be2d80",
  1218 => x"d19c08b2",
  1219 => x"3881ff0b",
  1220 => x"d40cd408",
  1221 => x"5381ff0b",
  1222 => x"d40c81ff",
  1223 => x"0bd40c81",
  1224 => x"ff0bd40c",
  1225 => x"81ff0bd4",
  1226 => x"0c72862a",
  1227 => x"70810676",
  1228 => x"56515372",
  1229 => x"963880d1",
  1230 => x"9c0854a6",
  1231 => x"cb047382",
  1232 => x"2efedb38",
  1233 => x"ff145473",
  1234 => x"fee73873",
  1235 => x"80d28c0c",
  1236 => x"738b3881",
  1237 => x"5287fc80",
  1238 => x"d051a2be",
  1239 => x"2d81ff0b",
  1240 => x"d40cd008",
  1241 => x"708f2a70",
  1242 => x"81065151",
  1243 => x"5372f338",
  1244 => x"72d00c81",
  1245 => x"ff0bd40c",
  1246 => x"81537280",
  1247 => x"d19c0c02",
  1248 => x"94050d04",
  1249 => x"02e8050d",
  1250 => x"78558056",
  1251 => x"81ff0bd4",
  1252 => x"0cd00870",
  1253 => x"8f2a7081",
  1254 => x"06515153",
  1255 => x"72f33882",
  1256 => x"810bd00c",
  1257 => x"81ff0bd4",
  1258 => x"0c775287",
  1259 => x"fc80d151",
  1260 => x"a2be2d80",
  1261 => x"dbc6df54",
  1262 => x"80d19c08",
  1263 => x"802e8b38",
  1264 => x"80c7f051",
  1265 => x"86c52da8",
  1266 => x"9e0481ff",
  1267 => x"0bd40cd4",
  1268 => x"087081ff",
  1269 => x"06515372",
  1270 => x"81fe2e09",
  1271 => x"81069e38",
  1272 => x"80ff53a1",
  1273 => x"ef2d80d1",
  1274 => x"9c087570",
  1275 => x"8405570c",
  1276 => x"ff135372",
  1277 => x"8025ec38",
  1278 => x"8156a883",
  1279 => x"04ff1454",
  1280 => x"73c83881",
  1281 => x"ff0bd40c",
  1282 => x"81ff0bd4",
  1283 => x"0cd00870",
  1284 => x"8f2a7081",
  1285 => x"06515153",
  1286 => x"72f33872",
  1287 => x"d00c7580",
  1288 => x"d19c0c02",
  1289 => x"98050d04",
  1290 => x"02e8050d",
  1291 => x"77797b58",
  1292 => x"55558053",
  1293 => x"727625a3",
  1294 => x"38747081",
  1295 => x"055680f5",
  1296 => x"2d747081",
  1297 => x"055680f5",
  1298 => x"2d525271",
  1299 => x"712e8638",
  1300 => x"8151a8dd",
  1301 => x"04811353",
  1302 => x"a8b40480",
  1303 => x"517080d1",
  1304 => x"9c0c0298",
  1305 => x"050d0402",
  1306 => x"ec050d76",
  1307 => x"5574802e",
  1308 => x"80c2389a",
  1309 => x"1580e02d",
  1310 => x"51b6fc2d",
  1311 => x"80d19c08",
  1312 => x"80d19c08",
  1313 => x"80d8c00c",
  1314 => x"80d19c08",
  1315 => x"545480d8",
  1316 => x"9c08802e",
  1317 => x"9a389415",
  1318 => x"80e02d51",
  1319 => x"b6fc2d80",
  1320 => x"d19c0890",
  1321 => x"2b83fff0",
  1322 => x"0a067075",
  1323 => x"07515372",
  1324 => x"80d8c00c",
  1325 => x"80d8c008",
  1326 => x"5372802e",
  1327 => x"9d3880d8",
  1328 => x"9408fe14",
  1329 => x"712980d8",
  1330 => x"a8080580",
  1331 => x"d8c40c70",
  1332 => x"842b80d8",
  1333 => x"a00c54aa",
  1334 => x"880480d8",
  1335 => x"ac0880d8",
  1336 => x"c00c80d8",
  1337 => x"b00880d8",
  1338 => x"c40c80d8",
  1339 => x"9c08802e",
  1340 => x"8b3880d8",
  1341 => x"9408842b",
  1342 => x"53aa8304",
  1343 => x"80d8b408",
  1344 => x"842b5372",
  1345 => x"80d8a00c",
  1346 => x"0294050d",
  1347 => x"0402d805",
  1348 => x"0d800b80",
  1349 => x"d89c0c84",
  1350 => x"54a4822d",
  1351 => x"80d19c08",
  1352 => x"802e9738",
  1353 => x"80d29052",
  1354 => x"8051a784",
  1355 => x"2d80d19c",
  1356 => x"08802e86",
  1357 => x"38fe54aa",
  1358 => x"c204ff14",
  1359 => x"54738024",
  1360 => x"d838738d",
  1361 => x"3880c880",
  1362 => x"5186c52d",
  1363 => x"7355b097",
  1364 => x"04805681",
  1365 => x"0b80d8c8",
  1366 => x"0c885380",
  1367 => x"c8945280",
  1368 => x"d2c651a8",
  1369 => x"a82d80d1",
  1370 => x"9c08762e",
  1371 => x"09810689",
  1372 => x"3880d19c",
  1373 => x"0880d8c8",
  1374 => x"0c885380",
  1375 => x"c8a05280",
  1376 => x"d2e251a8",
  1377 => x"a82d80d1",
  1378 => x"9c088938",
  1379 => x"80d19c08",
  1380 => x"80d8c80c",
  1381 => x"80d8c808",
  1382 => x"802e8181",
  1383 => x"3880d5d6",
  1384 => x"0b80f52d",
  1385 => x"80d5d70b",
  1386 => x"80f52d71",
  1387 => x"982b7190",
  1388 => x"2b0780d5",
  1389 => x"d80b80f5",
  1390 => x"2d70882b",
  1391 => x"720780d5",
  1392 => x"d90b80f5",
  1393 => x"2d710780",
  1394 => x"d68e0b80",
  1395 => x"f52d80d6",
  1396 => x"8f0b80f5",
  1397 => x"2d71882b",
  1398 => x"07535f54",
  1399 => x"525a5657",
  1400 => x"557381ab",
  1401 => x"aa2e0981",
  1402 => x"068e3875",
  1403 => x"51b6cb2d",
  1404 => x"80d19c08",
  1405 => x"56ac8604",
  1406 => x"7382d4d5",
  1407 => x"2e883880",
  1408 => x"c8ac51ac",
  1409 => x"d20480d2",
  1410 => x"90527551",
  1411 => x"a7842d80",
  1412 => x"d19c0855",
  1413 => x"80d19c08",
  1414 => x"802e83fb",
  1415 => x"38885380",
  1416 => x"c8a05280",
  1417 => x"d2e251a8",
  1418 => x"a82d80d1",
  1419 => x"9c088a38",
  1420 => x"810b80d8",
  1421 => x"9c0cacd8",
  1422 => x"04885380",
  1423 => x"c8945280",
  1424 => x"d2c651a8",
  1425 => x"a82d80d1",
  1426 => x"9c08802e",
  1427 => x"8b3880c8",
  1428 => x"c05186c5",
  1429 => x"2dadb704",
  1430 => x"80d68e0b",
  1431 => x"80f52d54",
  1432 => x"7380d52e",
  1433 => x"09810680",
  1434 => x"ce3880d6",
  1435 => x"8f0b80f5",
  1436 => x"2d547381",
  1437 => x"aa2e0981",
  1438 => x"06bd3880",
  1439 => x"0b80d290",
  1440 => x"0b80f52d",
  1441 => x"56547481",
  1442 => x"e92e8338",
  1443 => x"81547481",
  1444 => x"eb2e8c38",
  1445 => x"80557375",
  1446 => x"2e098106",
  1447 => x"82f93880",
  1448 => x"d29b0b80",
  1449 => x"f52d5574",
  1450 => x"8e3880d2",
  1451 => x"9c0b80f5",
  1452 => x"2d547382",
  1453 => x"2e863880",
  1454 => x"55b09704",
  1455 => x"80d29d0b",
  1456 => x"80f52d70",
  1457 => x"80d8940c",
  1458 => x"ff0580d8",
  1459 => x"980c80d2",
  1460 => x"9e0b80f5",
  1461 => x"2d80d29f",
  1462 => x"0b80f52d",
  1463 => x"58760577",
  1464 => x"82802905",
  1465 => x"7080d8a4",
  1466 => x"0c80d2a0",
  1467 => x"0b80f52d",
  1468 => x"7080d8b8",
  1469 => x"0c80d89c",
  1470 => x"08595758",
  1471 => x"76802e81",
  1472 => x"b7388853",
  1473 => x"80c8a052",
  1474 => x"80d2e251",
  1475 => x"a8a82d80",
  1476 => x"d19c0882",
  1477 => x"823880d8",
  1478 => x"94087084",
  1479 => x"2b80d8a0",
  1480 => x"0c7080d8",
  1481 => x"b40c80d2",
  1482 => x"b50b80f5",
  1483 => x"2d80d2b4",
  1484 => x"0b80f52d",
  1485 => x"71828029",
  1486 => x"0580d2b6",
  1487 => x"0b80f52d",
  1488 => x"70848080",
  1489 => x"291280d2",
  1490 => x"b70b80f5",
  1491 => x"2d708180",
  1492 => x"0a291270",
  1493 => x"80d8bc0c",
  1494 => x"80d8b808",
  1495 => x"712980d8",
  1496 => x"a4080570",
  1497 => x"80d8a80c",
  1498 => x"80d2bd0b",
  1499 => x"80f52d80",
  1500 => x"d2bc0b80",
  1501 => x"f52d7182",
  1502 => x"80290580",
  1503 => x"d2be0b80",
  1504 => x"f52d7084",
  1505 => x"80802912",
  1506 => x"80d2bf0b",
  1507 => x"80f52d70",
  1508 => x"982b81f0",
  1509 => x"0a067205",
  1510 => x"7080d8ac",
  1511 => x"0cfe117e",
  1512 => x"29770580",
  1513 => x"d8b00c52",
  1514 => x"59524354",
  1515 => x"5e515259",
  1516 => x"525d5759",
  1517 => x"57b09004",
  1518 => x"80d2a20b",
  1519 => x"80f52d80",
  1520 => x"d2a10b80",
  1521 => x"f52d7182",
  1522 => x"80290570",
  1523 => x"80d8a00c",
  1524 => x"70a02983",
  1525 => x"ff057089",
  1526 => x"2a7080d8",
  1527 => x"b40c80d2",
  1528 => x"a70b80f5",
  1529 => x"2d80d2a6",
  1530 => x"0b80f52d",
  1531 => x"71828029",
  1532 => x"057080d8",
  1533 => x"bc0c7b71",
  1534 => x"291e7080",
  1535 => x"d8b00c7d",
  1536 => x"80d8ac0c",
  1537 => x"730580d8",
  1538 => x"a80c555e",
  1539 => x"51515555",
  1540 => x"8051a8e7",
  1541 => x"2d815574",
  1542 => x"80d19c0c",
  1543 => x"02a8050d",
  1544 => x"0402ec05",
  1545 => x"0d767087",
  1546 => x"2c7180ff",
  1547 => x"06555654",
  1548 => x"80d89c08",
  1549 => x"8a387388",
  1550 => x"2c7481ff",
  1551 => x"06545580",
  1552 => x"d2905280",
  1553 => x"d8a40815",
  1554 => x"51a7842d",
  1555 => x"80d19c08",
  1556 => x"5480d19c",
  1557 => x"08802eb8",
  1558 => x"3880d89c",
  1559 => x"08802e9a",
  1560 => x"38728429",
  1561 => x"80d29005",
  1562 => x"70085253",
  1563 => x"b6cb2d80",
  1564 => x"d19c08f0",
  1565 => x"0a0653b1",
  1566 => x"8e047210",
  1567 => x"80d29005",
  1568 => x"7080e02d",
  1569 => x"5253b6fc",
  1570 => x"2d80d19c",
  1571 => x"08537254",
  1572 => x"7380d19c",
  1573 => x"0c029405",
  1574 => x"0d0402e0",
  1575 => x"050d7970",
  1576 => x"842c80d8",
  1577 => x"c4080571",
  1578 => x"8f065255",
  1579 => x"53728a38",
  1580 => x"80d29052",
  1581 => x"7351a784",
  1582 => x"2d72a029",
  1583 => x"80d29005",
  1584 => x"54807480",
  1585 => x"f52d5653",
  1586 => x"74732e83",
  1587 => x"38815374",
  1588 => x"81e52e81",
  1589 => x"f4388170",
  1590 => x"74065458",
  1591 => x"72802e81",
  1592 => x"e8388b14",
  1593 => x"80f52d70",
  1594 => x"832a7906",
  1595 => x"5856769b",
  1596 => x"3880cfe0",
  1597 => x"08537289",
  1598 => x"387280d6",
  1599 => x"900b81b7",
  1600 => x"2d7680cf",
  1601 => x"e00c7353",
  1602 => x"b3cb0475",
  1603 => x"8f2e0981",
  1604 => x"0681b638",
  1605 => x"749f068d",
  1606 => x"2980d683",
  1607 => x"11515381",
  1608 => x"1480f52d",
  1609 => x"73708105",
  1610 => x"5581b72d",
  1611 => x"831480f5",
  1612 => x"2d737081",
  1613 => x"055581b7",
  1614 => x"2d851480",
  1615 => x"f52d7370",
  1616 => x"81055581",
  1617 => x"b72d8714",
  1618 => x"80f52d73",
  1619 => x"70810555",
  1620 => x"81b72d89",
  1621 => x"1480f52d",
  1622 => x"73708105",
  1623 => x"5581b72d",
  1624 => x"8e1480f5",
  1625 => x"2d737081",
  1626 => x"055581b7",
  1627 => x"2d901480",
  1628 => x"f52d7370",
  1629 => x"81055581",
  1630 => x"b72d9214",
  1631 => x"80f52d73",
  1632 => x"70810555",
  1633 => x"81b72d94",
  1634 => x"1480f52d",
  1635 => x"73708105",
  1636 => x"5581b72d",
  1637 => x"961480f5",
  1638 => x"2d737081",
  1639 => x"055581b7",
  1640 => x"2d981480",
  1641 => x"f52d7370",
  1642 => x"81055581",
  1643 => x"b72d9c14",
  1644 => x"80f52d73",
  1645 => x"70810555",
  1646 => x"81b72d9e",
  1647 => x"1480f52d",
  1648 => x"7381b72d",
  1649 => x"7780cfe0",
  1650 => x"0c805372",
  1651 => x"80d19c0c",
  1652 => x"02a0050d",
  1653 => x"0402cc05",
  1654 => x"0d7e605e",
  1655 => x"5a800b80",
  1656 => x"d8c00880",
  1657 => x"d8c40859",
  1658 => x"5c568058",
  1659 => x"80d8a008",
  1660 => x"782e81b8",
  1661 => x"38778f06",
  1662 => x"a0175754",
  1663 => x"73913880",
  1664 => x"d2905276",
  1665 => x"51811757",
  1666 => x"a7842d80",
  1667 => x"d2905680",
  1668 => x"7680f52d",
  1669 => x"56547474",
  1670 => x"2e833881",
  1671 => x"547481e5",
  1672 => x"2e80fd38",
  1673 => x"81707506",
  1674 => x"555c7380",
  1675 => x"2e80f138",
  1676 => x"8b1680f5",
  1677 => x"2d980659",
  1678 => x"7880e538",
  1679 => x"8b537c52",
  1680 => x"7551a8a8",
  1681 => x"2d80d19c",
  1682 => x"0880d538",
  1683 => x"9c160851",
  1684 => x"b6cb2d80",
  1685 => x"d19c0884",
  1686 => x"1b0c9a16",
  1687 => x"80e02d51",
  1688 => x"b6fc2d80",
  1689 => x"d19c0880",
  1690 => x"d19c0888",
  1691 => x"1c0c80d1",
  1692 => x"9c085555",
  1693 => x"80d89c08",
  1694 => x"802e9938",
  1695 => x"941680e0",
  1696 => x"2d51b6fc",
  1697 => x"2d80d19c",
  1698 => x"08902b83",
  1699 => x"fff00a06",
  1700 => x"70165154",
  1701 => x"73881b0c",
  1702 => x"787a0c7b",
  1703 => x"54b5e804",
  1704 => x"81185880",
  1705 => x"d8a00878",
  1706 => x"26feca38",
  1707 => x"80d89c08",
  1708 => x"802eb338",
  1709 => x"7a51b0a1",
  1710 => x"2d80d19c",
  1711 => x"0880d19c",
  1712 => x"0880ffff",
  1713 => x"fff80655",
  1714 => x"5b7380ff",
  1715 => x"fffff82e",
  1716 => x"953880d1",
  1717 => x"9c08fe05",
  1718 => x"80d89408",
  1719 => x"2980d8a8",
  1720 => x"080557b3",
  1721 => x"ea048054",
  1722 => x"7380d19c",
  1723 => x"0c02b405",
  1724 => x"0d0402f4",
  1725 => x"050d7470",
  1726 => x"08810571",
  1727 => x"0c700880",
  1728 => x"d8980806",
  1729 => x"5353718f",
  1730 => x"38881308",
  1731 => x"51b0a12d",
  1732 => x"80d19c08",
  1733 => x"88140c81",
  1734 => x"0b80d19c",
  1735 => x"0c028c05",
  1736 => x"0d0402f0",
  1737 => x"050d7588",
  1738 => x"1108fe05",
  1739 => x"80d89408",
  1740 => x"2980d8a8",
  1741 => x"08117208",
  1742 => x"80d89808",
  1743 => x"06057955",
  1744 => x"535454a7",
  1745 => x"842d0290",
  1746 => x"050d0402",
  1747 => x"f4050d74",
  1748 => x"70882a83",
  1749 => x"fe800670",
  1750 => x"72982a07",
  1751 => x"72882b87",
  1752 => x"fc808006",
  1753 => x"73982b81",
  1754 => x"f00a0671",
  1755 => x"73070780",
  1756 => x"d19c0c56",
  1757 => x"51535102",
  1758 => x"8c050d04",
  1759 => x"02f8050d",
  1760 => x"028e0580",
  1761 => x"f52d7488",
  1762 => x"2b077083",
  1763 => x"ffff0680",
  1764 => x"d19c0c51",
  1765 => x"0288050d",
  1766 => x"0402f405",
  1767 => x"0d747678",
  1768 => x"53545280",
  1769 => x"71259738",
  1770 => x"72708105",
  1771 => x"5480f52d",
  1772 => x"72708105",
  1773 => x"5481b72d",
  1774 => x"ff115170",
  1775 => x"eb388072",
  1776 => x"81b72d02",
  1777 => x"8c050d04",
  1778 => x"02e8050d",
  1779 => x"77568070",
  1780 => x"56547376",
  1781 => x"24b63880",
  1782 => x"d8a00874",
  1783 => x"2eae3873",
  1784 => x"51b19a2d",
  1785 => x"80d19c08",
  1786 => x"80d19c08",
  1787 => x"09810570",
  1788 => x"80d19c08",
  1789 => x"079f2a77",
  1790 => x"05811757",
  1791 => x"57535374",
  1792 => x"76248938",
  1793 => x"80d8a008",
  1794 => x"7426d438",
  1795 => x"7280d19c",
  1796 => x"0c029805",
  1797 => x"0d0402ec",
  1798 => x"050d80d1",
  1799 => x"98081751",
  1800 => x"b7c82d80",
  1801 => x"d19c0855",
  1802 => x"80d19c08",
  1803 => x"802ea238",
  1804 => x"8b5380d1",
  1805 => x"9c085280",
  1806 => x"d69051b7",
  1807 => x"992d80d8",
  1808 => x"cc085473",
  1809 => x"802e8a38",
  1810 => x"88155280",
  1811 => x"d6905173",
  1812 => x"2d029405",
  1813 => x"0d0402dc",
  1814 => x"050d8070",
  1815 => x"5a557480",
  1816 => x"d1980825",
  1817 => x"b43880d8",
  1818 => x"a008752e",
  1819 => x"ac387851",
  1820 => x"b19a2d80",
  1821 => x"d19c0809",
  1822 => x"81057080",
  1823 => x"d19c0807",
  1824 => x"9f2a7605",
  1825 => x"811b5b56",
  1826 => x"547480d1",
  1827 => x"98082589",
  1828 => x"3880d8a0",
  1829 => x"087926d6",
  1830 => x"38805578",
  1831 => x"80d8a008",
  1832 => x"2781db38",
  1833 => x"7851b19a",
  1834 => x"2d80d19c",
  1835 => x"08802e81",
  1836 => x"ad3880d1",
  1837 => x"9c088b05",
  1838 => x"80f52d70",
  1839 => x"842a7081",
  1840 => x"06771078",
  1841 => x"842b80d6",
  1842 => x"900b80f5",
  1843 => x"2d5c5c53",
  1844 => x"51555673",
  1845 => x"802e80cb",
  1846 => x"38741682",
  1847 => x"2bbba20b",
  1848 => x"80cfec12",
  1849 => x"0c547775",
  1850 => x"311080d8",
  1851 => x"d0115556",
  1852 => x"90747081",
  1853 => x"055681b7",
  1854 => x"2da07481",
  1855 => x"b72d7681",
  1856 => x"ff068116",
  1857 => x"58547380",
  1858 => x"2e8a389c",
  1859 => x"5380d690",
  1860 => x"52ba9b04",
  1861 => x"8b5380d1",
  1862 => x"9c085280",
  1863 => x"d8d21651",
  1864 => x"bad60474",
  1865 => x"16822bb8",
  1866 => x"960b80cf",
  1867 => x"ec120c54",
  1868 => x"7681ff06",
  1869 => x"81165854",
  1870 => x"73802e8a",
  1871 => x"389c5380",
  1872 => x"d69052ba",
  1873 => x"cd048b53",
  1874 => x"80d19c08",
  1875 => x"52777531",
  1876 => x"1080d8d0",
  1877 => x"05517655",
  1878 => x"b7992dba",
  1879 => x"f3047490",
  1880 => x"29753170",
  1881 => x"1080d8d0",
  1882 => x"05515480",
  1883 => x"d19c0874",
  1884 => x"81b72d81",
  1885 => x"1959748b",
  1886 => x"24a338b9",
  1887 => x"9b047490",
  1888 => x"29753170",
  1889 => x"1080d8d0",
  1890 => x"058c7731",
  1891 => x"57515480",
  1892 => x"7481b72d",
  1893 => x"9e14ff16",
  1894 => x"565474f3",
  1895 => x"3802a405",
  1896 => x"0d0402fc",
  1897 => x"050d80d1",
  1898 => x"98081351",
  1899 => x"b7c82d80",
  1900 => x"d19c0880",
  1901 => x"2e893880",
  1902 => x"d19c0851",
  1903 => x"a8e72d80",
  1904 => x"0b80d198",
  1905 => x"0cb8d62d",
  1906 => x"93b82d02",
  1907 => x"84050d04",
  1908 => x"02fc050d",
  1909 => x"725170fd",
  1910 => x"2eb03870",
  1911 => x"fd248a38",
  1912 => x"70fc2e80",
  1913 => x"cc38bcbb",
  1914 => x"0470fe2e",
  1915 => x"b73870ff",
  1916 => x"2e098106",
  1917 => x"80c53880",
  1918 => x"d1980851",
  1919 => x"70802ebb",
  1920 => x"38ff1180",
  1921 => x"d1980cbc",
  1922 => x"bb0480d1",
  1923 => x"9808f405",
  1924 => x"7080d198",
  1925 => x"0c517080",
  1926 => x"25a13880",
  1927 => x"0b80d198",
  1928 => x"0cbcbb04",
  1929 => x"80d19808",
  1930 => x"810580d1",
  1931 => x"980cbcbb",
  1932 => x"0480d198",
  1933 => x"088c0580",
  1934 => x"d1980cb8",
  1935 => x"d62d93b8",
  1936 => x"2d028405",
  1937 => x"0d0402fc",
  1938 => x"050d800b",
  1939 => x"80d1980c",
  1940 => x"b8d62d92",
  1941 => x"a62d80d1",
  1942 => x"9c0880d1",
  1943 => x"880c80cf",
  1944 => x"e45194de",
  1945 => x"2d028405",
  1946 => x"0d0402fc",
  1947 => x"050d810b",
  1948 => x"80c8d80c",
  1949 => x"7251bcc6",
  1950 => x"2d028405",
  1951 => x"0d0402fc",
  1952 => x"050d800b",
  1953 => x"80c8d80c",
  1954 => x"7251bcc6",
  1955 => x"2d028405",
  1956 => x"0d047180",
  1957 => x"d8cc0c04",
  1958 => x"00ffffff",
  1959 => x"ff00ffff",
  1960 => x"ffff00ff",
  1961 => x"ffffff00",
  1962 => x"4b455953",
  1963 => x"50312020",
  1964 => x"20202000",
  1965 => x"00000000",
  1966 => x"4b455953",
  1967 => x"50322020",
  1968 => x"20202000",
  1969 => x"00000000",
  1970 => x"3d3d2056",
  1971 => x"6964656f",
  1972 => x"70616320",
  1973 => x"666f7220",
  1974 => x"5a58444f",
  1975 => x"53203d3d",
  1976 => x"00000000",
  1977 => x"3d3d3d3d",
  1978 => x"3d3d3d3d",
  1979 => x"3d3d3d3d",
  1980 => x"3d3d3d3d",
  1981 => x"3d3d3d3d",
  1982 => x"3d3d3d3d",
  1983 => x"00000000",
  1984 => x"52657365",
  1985 => x"74000000",
  1986 => x"5363616e",
  1987 => x"6c696e65",
  1988 => x"73000000",
  1989 => x"53776170",
  1990 => x"206a6f79",
  1991 => x"73746963",
  1992 => x"6b730000",
  1993 => x"4a6f696e",
  1994 => x"206a6f79",
  1995 => x"73746963",
  1996 => x"6b730000",
  1997 => x"4c6f6164",
  1998 => x"20636174",
  1999 => x"72696467",
  2000 => x"6520524f",
  2001 => x"4d201000",
  2002 => x"4c6f6164",
  2003 => x"20564443",
  2004 => x"20666f6e",
  2005 => x"74201000",
  2006 => x"48656c70",
  2007 => x"00000000",
  2008 => x"45786974",
  2009 => x"00000000",
  2010 => x"54686520",
  2011 => x"766f6963",
  2012 => x"653a204f",
  2013 => x"66660000",
  2014 => x"54686520",
  2015 => x"766f6963",
  2016 => x"653a204f",
  2017 => x"6e000000",
  2018 => x"436f6c6f",
  2019 => x"72206d6f",
  2020 => x"64653a20",
  2021 => x"436f6c6f",
  2022 => x"72000000",
  2023 => x"436f6c6f",
  2024 => x"72206d6f",
  2025 => x"64653a20",
  2026 => x"4d6f6e6f",
  2027 => x"6368726f",
  2028 => x"6d650000",
  2029 => x"436f6c6f",
  2030 => x"72206d6f",
  2031 => x"64653a20",
  2032 => x"47726565",
  2033 => x"6e207068",
  2034 => x"6f737068",
  2035 => x"6f720000",
  2036 => x"436f6c6f",
  2037 => x"72206d6f",
  2038 => x"64653a20",
  2039 => x"416d6265",
  2040 => x"72206d6f",
  2041 => x"6e6f6368",
  2042 => x"726f6d65",
  2043 => x"00000000",
  2044 => x"4d6f6465",
  2045 => x"3a204f64",
  2046 => x"79737365",
  2047 => x"79322028",
  2048 => x"4e545343",
  2049 => x"29000000",
  2050 => x"4d6f6465",
  2051 => x"3a205669",
  2052 => x"64656f70",
  2053 => x"61632028",
  2054 => x"50414c29",
  2055 => x"00000000",
  2056 => x"3d3d2056",
  2057 => x"6964656f",
  2058 => x"70616320",
  2059 => x"666f7220",
  2060 => x"5a58554e",
  2061 => x"4f203d3d",
  2062 => x"00000000",
  2063 => x"5a58554e",
  2064 => x"4f3a2073",
  2065 => x"696e676c",
  2066 => x"65206a6f",
  2067 => x"79737469",
  2068 => x"636b0000",
  2069 => x"5a58554e",
  2070 => x"4f3a2032",
  2071 => x"206a6f79",
  2072 => x"73746963",
  2073 => x"6b207370",
  2074 => x"6c697474",
  2075 => x"65720000",
  2076 => x"5a58554e",
  2077 => x"4f3a2032",
  2078 => x"206a6f79",
  2079 => x"73746963",
  2080 => x"6b205647",
  2081 => x"41324d00",
  2082 => x"524f4d20",
  2083 => x"6c6f6164",
  2084 => x"696e6720",
  2085 => x"6661696c",
  2086 => x"65640000",
  2087 => x"4f4b0000",
  2088 => x"3d3d3d20",
  2089 => x"56696465",
  2090 => x"6f706163",
  2091 => x"20537065",
  2092 => x"6369616c",
  2093 => x"2048454c",
  2094 => x"50203d3d",
  2095 => x"3d000000",
  2096 => x"3d3d3d3d",
  2097 => x"3d3d3d3d",
  2098 => x"3d3d3d3d",
  2099 => x"3d3d3d3d",
  2100 => x"3d3d3d3d",
  2101 => x"3d3d3d3d",
  2102 => x"3d3d3d3d",
  2103 => x"3d3d0000",
  2104 => x"5363726f",
  2105 => x"6c6c204c",
  2106 => x"6f636b3a",
  2107 => x"20636861",
  2108 => x"6e676520",
  2109 => x"62657477",
  2110 => x"65656e00",
  2111 => x"52474220",
  2112 => x"616e6420",
  2113 => x"56474120",
  2114 => x"76696465",
  2115 => x"6f206d6f",
  2116 => x"64650000",
  2117 => x"46333a20",
  2118 => x"536f6674",
  2119 => x"20526573",
  2120 => x"65740000",
  2121 => x"4374726c",
  2122 => x"2b416c74",
  2123 => x"2b426163",
  2124 => x"6b737061",
  2125 => x"63653a20",
  2126 => x"48617264",
  2127 => x"20726573",
  2128 => x"65740000",
  2129 => x"45736320",
  2130 => x"6f72206a",
  2131 => x"6f797374",
  2132 => x"69636b20",
  2133 => x"62742e32",
  2134 => x"3a20746f",
  2135 => x"2073686f",
  2136 => x"77000000",
  2137 => x"6f722068",
  2138 => x"69646520",
  2139 => x"74686520",
  2140 => x"6f707469",
  2141 => x"6f6e7320",
  2142 => x"6d656e75",
  2143 => x"2e000000",
  2144 => x"57415344",
  2145 => x"202f2063",
  2146 => x"7572736f",
  2147 => x"72206b65",
  2148 => x"7973202f",
  2149 => x"206a6f79",
  2150 => x"73746963",
  2151 => x"6b000000",
  2152 => x"746f2073",
  2153 => x"656c6563",
  2154 => x"74206d65",
  2155 => x"6e75206f",
  2156 => x"7074696f",
  2157 => x"6e2e0000",
  2158 => x"456e7465",
  2159 => x"72202f20",
  2160 => x"46697265",
  2161 => x"20746f20",
  2162 => x"63686f6f",
  2163 => x"7365206f",
  2164 => x"7074696f",
  2165 => x"6e2e0000",
  2166 => x"496e206d",
  2167 => x"6f737420",
  2168 => x"67616d65",
  2169 => x"73207072",
  2170 => x"65737320",
  2171 => x"302d3920",
  2172 => x"61667465",
  2173 => x"72000000",
  2174 => x"6c6f6164",
  2175 => x"696e6720",
  2176 => x"6120524f",
  2177 => x"4d20746f",
  2178 => x"20706c61",
  2179 => x"79207468",
  2180 => x"65206761",
  2181 => x"6d650000",
  2182 => x"3d3d3d20",
  2183 => x"56696465",
  2184 => x"6f706163",
  2185 => x"20436f72",
  2186 => x"65204372",
  2187 => x"65646974",
  2188 => x"73203d3d",
  2189 => x"3d000000",
  2190 => x"3d3d3d3d",
  2191 => x"3d3d3d3d",
  2192 => x"3d3d3d3d",
  2193 => x"3d3d3d3d",
  2194 => x"3d3d3d3d",
  2195 => x"3d3d3d3d",
  2196 => x"3d3d3d3d",
  2197 => x"3d000000",
  2198 => x"5068696c",
  2199 => x"69707320",
  2200 => x"56696465",
  2201 => x"6f706163",
  2202 => x"202f204d",
  2203 => x"61676e61",
  2204 => x"766f7800",
  2205 => x"4f647973",
  2206 => x"73657932",
  2207 => x"20636f72",
  2208 => x"6520666f",
  2209 => x"72205a58",
  2210 => x"554e4f2c",
  2211 => x"205a5844",
  2212 => x"4f530000",
  2213 => x"616e6420",
  2214 => x"5a58444f",
  2215 => x"532b2062",
  2216 => x"6f617264",
  2217 => x"732e0000",
  2218 => x"4f726967",
  2219 => x"696e616c",
  2220 => x"20636f72",
  2221 => x"65206279",
  2222 => x"3a41726e",
  2223 => x"696d204c",
  2224 => x"61657567",
  2225 => x"65720000",
  2226 => x"506f7274",
  2227 => x"206d6164",
  2228 => x"65206279",
  2229 => x"3a20796f",
  2230 => x"6d626f70",
  2231 => x"72696d65",
  2232 => x"2c200000",
  2233 => x"2072616d",
  2234 => x"70613036",
  2235 => x"392c206e",
  2236 => x"6575726f",
  2237 => x"72756c65",
  2238 => x"7a2c2041",
  2239 => x"6e746f6e",
  2240 => x"696f0000",
  2241 => x"2053616e",
  2242 => x"6368657a",
  2243 => x"2c204176",
  2244 => x"6c697841",
  2245 => x"2c204d65",
  2246 => x"6a696173",
  2247 => x"33442c20",
  2248 => x"00000000",
  2249 => x"2057696c",
  2250 => x"636f3230",
  2251 => x"30392061",
  2252 => x"6e642042",
  2253 => x"656e6974",
  2254 => x"6f737300",
  2255 => x"53706563",
  2256 => x"69616c20",
  2257 => x"5468616e",
  2258 => x"6b732074",
  2259 => x"6f3a2052",
  2260 => x"656e6520",
  2261 => x"76616e20",
  2262 => x"00000000",
  2263 => x"2064656e",
  2264 => x"20456e64",
  2265 => x"656e2066",
  2266 => x"6f722068",
  2267 => x"69732069",
  2268 => x"6e666f20",
  2269 => x"6f6e2000",
  2270 => x"20766964",
  2271 => x"656f7061",
  2272 => x"632e6e6c",
  2273 => x"00000000",
  2274 => x"496e6974",
  2275 => x"69616c69",
  2276 => x"7a696e67",
  2277 => x"20534420",
  2278 => x"63617264",
  2279 => x"0a000000",
  2280 => x"16200000",
  2281 => x"14200000",
  2282 => x"15200000",
  2283 => x"53442069",
  2284 => x"6e69742e",
  2285 => x"2e2e0a00",
  2286 => x"53442063",
  2287 => x"61726420",
  2288 => x"72657365",
  2289 => x"74206661",
  2290 => x"696c6564",
  2291 => x"210a0000",
  2292 => x"53444843",
  2293 => x"20657272",
  2294 => x"6f72210a",
  2295 => x"00000000",
  2296 => x"57726974",
  2297 => x"65206661",
  2298 => x"696c6564",
  2299 => x"0a000000",
  2300 => x"52656164",
  2301 => x"20666169",
  2302 => x"6c65640a",
  2303 => x"00000000",
  2304 => x"43617264",
  2305 => x"20696e69",
  2306 => x"74206661",
  2307 => x"696c6564",
  2308 => x"0a000000",
  2309 => x"46415431",
  2310 => x"36202020",
  2311 => x"00000000",
  2312 => x"46415433",
  2313 => x"32202020",
  2314 => x"00000000",
  2315 => x"4e6f2070",
  2316 => x"61727469",
  2317 => x"74696f6e",
  2318 => x"20736967",
  2319 => x"0a000000",
  2320 => x"42616420",
  2321 => x"70617274",
  2322 => x"0a000000",
  2323 => x"4261636b",
  2324 => x"00000000",
  2325 => x"00000002",
  2326 => x"00000000",
  2327 => x"00000010",
  2328 => x"00000002",
  2329 => x"00001ec8",
  2330 => x"000003ab",
  2331 => x"00000002",
  2332 => x"00001ee4",
  2333 => x"000003ab",
  2334 => x"00000002",
  2335 => x"00001f00",
  2336 => x"0000037f",
  2337 => x"00000001",
  2338 => x"00001f08",
  2339 => x"00000000",
  2340 => x"00000001",
  2341 => x"00001f14",
  2342 => x"00000001",
  2343 => x"00000001",
  2344 => x"00001f24",
  2345 => x"00000002",
  2346 => x"00000002",
  2347 => x"00001f34",
  2348 => x"00001e7e",
  2349 => x"00000002",
  2350 => x"00001f48",
  2351 => x"00001e6a",
  2352 => x"00000003",
  2353 => x"00002520",
  2354 => x"00000002",
  2355 => x"00000003",
  2356 => x"00002510",
  2357 => x"00000004",
  2358 => x"00000003",
  2359 => x"00002508",
  2360 => x"00000002",
  2361 => x"00000002",
  2362 => x"00001f58",
  2363 => x"000003c6",
  2364 => x"00000002",
  2365 => x"00001f60",
  2366 => x"00000943",
  2367 => x"00000000",
  2368 => x"00000000",
  2369 => x"00000000",
  2370 => x"00001f68",
  2371 => x"00001f78",
  2372 => x"00001f88",
  2373 => x"00001f9c",
  2374 => x"00001fb4",
  2375 => x"00001fd0",
  2376 => x"00001ff0",
  2377 => x"00002008",
  2378 => x"00000002",
  2379 => x"00002020",
  2380 => x"000003ab",
  2381 => x"00000002",
  2382 => x"00001ee4",
  2383 => x"000003ab",
  2384 => x"00000002",
  2385 => x"00001f00",
  2386 => x"0000037f",
  2387 => x"00000001",
  2388 => x"00001f08",
  2389 => x"00000000",
  2390 => x"00000001",
  2391 => x"00001f14",
  2392 => x"00000001",
  2393 => x"00000001",
  2394 => x"00001f24",
  2395 => x"00000002",
  2396 => x"00000002",
  2397 => x"00001f34",
  2398 => x"00001e7e",
  2399 => x"00000002",
  2400 => x"00001f48",
  2401 => x"00001e6a",
  2402 => x"00000003",
  2403 => x"00002520",
  2404 => x"00000002",
  2405 => x"00000003",
  2406 => x"00002510",
  2407 => x"00000004",
  2408 => x"00000003",
  2409 => x"000025d0",
  2410 => x"00000003",
  2411 => x"00000002",
  2412 => x"00001f58",
  2413 => x"000003c6",
  2414 => x"00000002",
  2415 => x"00001f60",
  2416 => x"00000943",
  2417 => x"00000000",
  2418 => x"00000000",
  2419 => x"00000000",
  2420 => x"0000203c",
  2421 => x"00002054",
  2422 => x"00002070",
  2423 => x"00000004",
  2424 => x"00002088",
  2425 => x"000025dc",
  2426 => x"00000004",
  2427 => x"0000209c",
  2428 => x"000028c4",
  2429 => x"00000000",
  2430 => x"00000000",
  2431 => x"00000000",
  2432 => x"00000002",
  2433 => x"000020a0",
  2434 => x"000003aa",
  2435 => x"00000002",
  2436 => x"000020c0",
  2437 => x"000003aa",
  2438 => x"00000002",
  2439 => x"000020e0",
  2440 => x"000003aa",
  2441 => x"00000002",
  2442 => x"000020fc",
  2443 => x"000003aa",
  2444 => x"00000002",
  2445 => x"00002114",
  2446 => x"000003aa",
  2447 => x"00000002",
  2448 => x"00002124",
  2449 => x"000003aa",
  2450 => x"00000002",
  2451 => x"00002144",
  2452 => x"000003aa",
  2453 => x"00000002",
  2454 => x"00002164",
  2455 => x"000003aa",
  2456 => x"00000002",
  2457 => x"00002180",
  2458 => x"000003aa",
  2459 => x"00000002",
  2460 => x"000021a0",
  2461 => x"000003aa",
  2462 => x"00000002",
  2463 => x"000021b8",
  2464 => x"000003aa",
  2465 => x"00000002",
  2466 => x"000021d8",
  2467 => x"000003aa",
  2468 => x"00000002",
  2469 => x"000021f8",
  2470 => x"000003aa",
  2471 => x"00000004",
  2472 => x"0000209c",
  2473 => x"000028c4",
  2474 => x"00000000",
  2475 => x"00000000",
  2476 => x"00000000",
  2477 => x"00000002",
  2478 => x"00002218",
  2479 => x"000003aa",
  2480 => x"00000002",
  2481 => x"00002238",
  2482 => x"000003aa",
  2483 => x"00000002",
  2484 => x"00002258",
  2485 => x"000003aa",
  2486 => x"00000002",
  2487 => x"00002274",
  2488 => x"000003aa",
  2489 => x"00000002",
  2490 => x"00002294",
  2491 => x"000003aa",
  2492 => x"00000002",
  2493 => x"000022a8",
  2494 => x"000003aa",
  2495 => x"00000002",
  2496 => x"000022c8",
  2497 => x"000003aa",
  2498 => x"00000002",
  2499 => x"000022e4",
  2500 => x"000003aa",
  2501 => x"00000002",
  2502 => x"00002304",
  2503 => x"000003aa",
  2504 => x"00000002",
  2505 => x"00002324",
  2506 => x"000003aa",
  2507 => x"00000002",
  2508 => x"0000233c",
  2509 => x"000003aa",
  2510 => x"00000002",
  2511 => x"0000235c",
  2512 => x"000003aa",
  2513 => x"00000002",
  2514 => x"00002378",
  2515 => x"000003aa",
  2516 => x"00000004",
  2517 => x"0000209c",
  2518 => x"000028c4",
  2519 => x"00000000",
  2520 => x"00000000",
  2521 => x"00000000",
  2522 => x"00000000",
  2523 => x"00000000",
  2524 => x"00000000",
  2525 => x"00000000",
  2526 => x"00000000",
  2527 => x"00000000",
  2528 => x"00000000",
  2529 => x"00000000",
  2530 => x"00000000",
  2531 => x"00000000",
  2532 => x"00000000",
  2533 => x"00000000",
  2534 => x"00000000",
  2535 => x"00000000",
  2536 => x"00000000",
  2537 => x"00000000",
  2538 => x"00000000",
  2539 => x"00000000",
  2540 => x"00000006",
  2541 => x"00000043",
  2542 => x"00000042",
  2543 => x"0000003b",
  2544 => x"0000004b",
  2545 => x"00000033",
  2546 => x"0000001d",
  2547 => x"0000001b",
  2548 => x"0000001c",
  2549 => x"00000023",
  2550 => x"0000002b",
  2551 => x"00000000",
  2552 => x"00000000",
  2553 => x"00000002",
  2554 => x"00002c50",
  2555 => x"00001c16",
  2556 => x"00000002",
  2557 => x"00002c6e",
  2558 => x"00001c16",
  2559 => x"00000002",
  2560 => x"00002c8c",
  2561 => x"00001c16",
  2562 => x"00000002",
  2563 => x"00002caa",
  2564 => x"00001c16",
  2565 => x"00000002",
  2566 => x"00002cc8",
  2567 => x"00001c16",
  2568 => x"00000002",
  2569 => x"00002ce6",
  2570 => x"00001c16",
  2571 => x"00000002",
  2572 => x"00002d04",
  2573 => x"00001c16",
  2574 => x"00000002",
  2575 => x"00002d22",
  2576 => x"00001c16",
  2577 => x"00000002",
  2578 => x"00002d40",
  2579 => x"00001c16",
  2580 => x"00000002",
  2581 => x"00002d5e",
  2582 => x"00001c16",
  2583 => x"00000002",
  2584 => x"00002d7c",
  2585 => x"00001c16",
  2586 => x"00000002",
  2587 => x"00002d9a",
  2588 => x"00001c16",
  2589 => x"00000002",
  2590 => x"00002db8",
  2591 => x"00001c16",
  2592 => x"00000004",
  2593 => x"0000244c",
  2594 => x"00000000",
  2595 => x"00000000",
  2596 => x"00000000",
  2597 => x"00001dd0",
  2598 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

