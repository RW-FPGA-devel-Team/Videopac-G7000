-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb7",
     9 => x"a0080b0b",
    10 => x"0bb7a408",
    11 => x"0b0b0bb7",
    12 => x"a8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b7a80c0b",
    16 => x"0b0bb7a4",
    17 => x"0c0b0b0b",
    18 => x"b7a00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafb0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b7a07080",
    57 => x"c1d0278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e604",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb7b00c",
    65 => x"9f0bb7b4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b7b408ff",
    69 => x"05b7b40c",
    70 => x"b7b40880",
    71 => x"25eb38b7",
    72 => x"b008ff05",
    73 => x"b7b00cb7",
    74 => x"b0088025",
    75 => x"d738800b",
    76 => x"b7b40c80",
    77 => x"0bb7b00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb7b008",
    97 => x"258f3882",
    98 => x"bd2db7b0",
    99 => x"08ff05b7",
   100 => x"b00c82ff",
   101 => x"04b7b008",
   102 => x"b7b40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b7b008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b7b4",
   111 => x"088105b7",
   112 => x"b40cb7b4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb7b40c",
   116 => x"b7b00881",
   117 => x"05b7b00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b7",
   122 => x"b4088105",
   123 => x"b7b40cb7",
   124 => x"b408a02e",
   125 => x"0981068e",
   126 => x"38800bb7",
   127 => x"b40cb7b0",
   128 => x"088105b7",
   129 => x"b00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb7b8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb7b80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b7",
   169 => x"b8088407",
   170 => x"b7b80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb3a4",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b7b80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b7a00c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c8dcf2d",
   216 => x"0284050d",
   217 => x"0402fc05",
   218 => x"0dec5192",
   219 => x"710c86a4",
   220 => x"2d82710c",
   221 => x"0284050d",
   222 => x"0402d005",
   223 => x"0d7d5480",
   224 => x"5ba40bec",
   225 => x"0c7352b7",
   226 => x"bc51a6ee",
   227 => x"2db7a008",
   228 => x"7b2e81ab",
   229 => x"38b7c008",
   230 => x"70f80c89",
   231 => x"1580f52d",
   232 => x"8a1680f5",
   233 => x"2d718280",
   234 => x"29058817",
   235 => x"80f52d70",
   236 => x"84808029",
   237 => x"12f40c7e",
   238 => x"ff155c5e",
   239 => x"57555658",
   240 => x"767b2e8b",
   241 => x"38811a77",
   242 => x"812a585a",
   243 => x"76f738f7",
   244 => x"1a5a815b",
   245 => x"80782580",
   246 => x"e6387952",
   247 => x"7651848b",
   248 => x"2db88852",
   249 => x"b7bc51a9",
   250 => x"a42db7a0",
   251 => x"08802eb8",
   252 => x"38b8885c",
   253 => x"83fc597b",
   254 => x"7084055d",
   255 => x"087081ff",
   256 => x"0671882a",
   257 => x"7081ff06",
   258 => x"73902a70",
   259 => x"81ff0675",
   260 => x"982ae80c",
   261 => x"e80c58e8",
   262 => x"0c57e80c",
   263 => x"fc1a5a53",
   264 => x"788025d3",
   265 => x"3888af04",
   266 => x"b7a0085b",
   267 => x"848058b7",
   268 => x"bc51a8f7",
   269 => x"2dfc8018",
   270 => x"81185858",
   271 => x"87d40486",
   272 => x"b72d800b",
   273 => x"ec0c7a80",
   274 => x"2e8d38b3",
   275 => x"a8518fcc",
   276 => x"2d8dcf2d",
   277 => x"88dd04b4",
   278 => x"f0518fcc",
   279 => x"2d7ab7a0",
   280 => x"0c02b005",
   281 => x"0d0402ec",
   282 => x"050d850b",
   283 => x"ec0c8db0",
   284 => x"2d8a9a2d",
   285 => x"81f82d9e",
   286 => x"8b2db7a0",
   287 => x"08802e81",
   288 => x"843886f9",
   289 => x"51afab2d",
   290 => x"b3a8518f",
   291 => x"cc2d8dcf",
   292 => x"2d8aa62d",
   293 => x"8fdc2db3",
   294 => x"d40b80f5",
   295 => x"2d70892b",
   296 => x"8c8006b3",
   297 => x"e00b80f5",
   298 => x"2d70872b",
   299 => x"818006b3",
   300 => x"ec0b80f5",
   301 => x"2d701082",
   302 => x"06747307",
   303 => x"07b3f80b",
   304 => x"80f52d70",
   305 => x"852ba006",
   306 => x"b4840b80",
   307 => x"f52d708e",
   308 => x"2b818080",
   309 => x"06747307",
   310 => x"07b4900b",
   311 => x"80f52d70",
   312 => x"862b80c0",
   313 => x"067207fc",
   314 => x"0c535454",
   315 => x"54565452",
   316 => x"57575353",
   317 => x"8652b7a0",
   318 => x"088538b7",
   319 => x"a0085271",
   320 => x"ec0c8991",
   321 => x"04800bb7",
   322 => x"a00c0294",
   323 => x"050d0471",
   324 => x"980c04ff",
   325 => x"b008b7a0",
   326 => x"0c04810b",
   327 => x"ffb00c04",
   328 => x"800bffb0",
   329 => x"0c0402f4",
   330 => x"050d8ba8",
   331 => x"04b7a008",
   332 => x"81f02e09",
   333 => x"81068938",
   334 => x"810bb5d4",
   335 => x"0c8ba804",
   336 => x"b7a00881",
   337 => x"e02e0981",
   338 => x"06893881",
   339 => x"0bb5d80c",
   340 => x"8ba804b7",
   341 => x"a00852b5",
   342 => x"d808802e",
   343 => x"8838b7a0",
   344 => x"08818005",
   345 => x"5271842c",
   346 => x"728f0653",
   347 => x"53b5d408",
   348 => x"802e9938",
   349 => x"728429b5",
   350 => x"94057213",
   351 => x"81712b70",
   352 => x"09730806",
   353 => x"730c5153",
   354 => x"538b9e04",
   355 => x"728429b5",
   356 => x"94057213",
   357 => x"83712b72",
   358 => x"0807720c",
   359 => x"5353800b",
   360 => x"b5d80c80",
   361 => x"0bb5d40c",
   362 => x"b7c8518c",
   363 => x"a92db7a0",
   364 => x"08ff24fe",
   365 => x"f838800b",
   366 => x"b7a00c02",
   367 => x"8c050d04",
   368 => x"02f8050d",
   369 => x"b594528f",
   370 => x"51807270",
   371 => x"8405540c",
   372 => x"ff115170",
   373 => x"8025f238",
   374 => x"0288050d",
   375 => x"0402f005",
   376 => x"0d75518a",
   377 => x"a02d7082",
   378 => x"2cfc06b5",
   379 => x"94117210",
   380 => x"9e067108",
   381 => x"70722a70",
   382 => x"83068274",
   383 => x"2b700974",
   384 => x"06760c54",
   385 => x"51565753",
   386 => x"51538a9a",
   387 => x"2d71b7a0",
   388 => x"0c029005",
   389 => x"0d0402fc",
   390 => x"050d7251",
   391 => x"80710c80",
   392 => x"0b84120c",
   393 => x"0284050d",
   394 => x"0402f005",
   395 => x"0d757008",
   396 => x"84120853",
   397 => x"5353ff54",
   398 => x"71712ea8",
   399 => x"388aa02d",
   400 => x"84130870",
   401 => x"84291488",
   402 => x"11700870",
   403 => x"81ff0684",
   404 => x"18088111",
   405 => x"8706841a",
   406 => x"0c535155",
   407 => x"5151518a",
   408 => x"9a2d7154",
   409 => x"73b7a00c",
   410 => x"0290050d",
   411 => x"0402f805",
   412 => x"0d8aa02d",
   413 => x"e008708b",
   414 => x"2a708106",
   415 => x"51525270",
   416 => x"802e9d38",
   417 => x"b7c80870",
   418 => x"8429b7d0",
   419 => x"057381ff",
   420 => x"06710c51",
   421 => x"51b7c808",
   422 => x"81118706",
   423 => x"b7c80c51",
   424 => x"800bb7f0",
   425 => x"0c8a932d",
   426 => x"8a9a2d02",
   427 => x"88050d04",
   428 => x"02fc050d",
   429 => x"b7c8518c",
   430 => x"962d8bc0",
   431 => x"2d8ced51",
   432 => x"8a8f2d02",
   433 => x"84050d04",
   434 => x"b7f408b7",
   435 => x"a00c0402",
   436 => x"fc050d8d",
   437 => x"d9048aa6",
   438 => x"2d80f651",
   439 => x"8bdd2db7",
   440 => x"a008f338",
   441 => x"80da518b",
   442 => x"dd2db7a0",
   443 => x"08e838b7",
   444 => x"a008b5e0",
   445 => x"0cb7a008",
   446 => x"5184f02d",
   447 => x"0284050d",
   448 => x"0402ec05",
   449 => x"0d765480",
   450 => x"52870b88",
   451 => x"1580f52d",
   452 => x"56537472",
   453 => x"248338a0",
   454 => x"53725182",
   455 => x"f92d8112",
   456 => x"8b1580f5",
   457 => x"2d545272",
   458 => x"7225de38",
   459 => x"0294050d",
   460 => x"0402f005",
   461 => x"0db7f408",
   462 => x"5481f82d",
   463 => x"800bb7f8",
   464 => x"0c730880",
   465 => x"2e818038",
   466 => x"820bb7b4",
   467 => x"0cb7f808",
   468 => x"8f06b7b0",
   469 => x"0c730852",
   470 => x"71832e96",
   471 => x"38718326",
   472 => x"89387181",
   473 => x"2eaf388f",
   474 => x"b2047185",
   475 => x"2e9f388f",
   476 => x"b2048814",
   477 => x"80f52d84",
   478 => x"1508b1f0",
   479 => x"53545285",
   480 => x"fe2d7184",
   481 => x"29137008",
   482 => x"52528fb6",
   483 => x"0473518e",
   484 => x"812d8fb2",
   485 => x"04b5dc08",
   486 => x"8815082c",
   487 => x"70810651",
   488 => x"5271802e",
   489 => x"8738b1f4",
   490 => x"518faf04",
   491 => x"b1f85185",
   492 => x"fe2d8414",
   493 => x"085185fe",
   494 => x"2db7f808",
   495 => x"8105b7f8",
   496 => x"0c8c1454",
   497 => x"8ec10402",
   498 => x"90050d04",
   499 => x"71b7f40c",
   500 => x"8eb12db7",
   501 => x"f808ff05",
   502 => x"b7fc0c04",
   503 => x"02e8050d",
   504 => x"b7f408b8",
   505 => x"80085755",
   506 => x"87518bdd",
   507 => x"2db7a008",
   508 => x"812a7081",
   509 => x"06515271",
   510 => x"802ea038",
   511 => x"9082048a",
   512 => x"a62d8751",
   513 => x"8bdd2db7",
   514 => x"a008f438",
   515 => x"b5e00881",
   516 => x"3270b5e0",
   517 => x"0c705252",
   518 => x"84f02d80",
   519 => x"fe518bdd",
   520 => x"2db7a008",
   521 => x"802ea638",
   522 => x"b5e00880",
   523 => x"2e913880",
   524 => x"0bb5e00c",
   525 => x"805184f0",
   526 => x"2d90bf04",
   527 => x"8aa62d80",
   528 => x"fe518bdd",
   529 => x"2db7a008",
   530 => x"f33886e5",
   531 => x"2db5e008",
   532 => x"903881fd",
   533 => x"518bdd2d",
   534 => x"81fa518b",
   535 => x"dd2d9692",
   536 => x"0481f551",
   537 => x"8bdd2db7",
   538 => x"a008812a",
   539 => x"70810651",
   540 => x"5271802e",
   541 => x"af38b7fc",
   542 => x"08527180",
   543 => x"2e8938ff",
   544 => x"12b7fc0c",
   545 => x"91a404b7",
   546 => x"f80810b7",
   547 => x"f8080570",
   548 => x"84291651",
   549 => x"52881208",
   550 => x"802e8938",
   551 => x"ff518812",
   552 => x"0852712d",
   553 => x"81f2518b",
   554 => x"dd2db7a0",
   555 => x"08812a70",
   556 => x"81065152",
   557 => x"71802eb1",
   558 => x"38b7f808",
   559 => x"ff11b7fc",
   560 => x"08565353",
   561 => x"73722589",
   562 => x"388114b7",
   563 => x"fc0c91e9",
   564 => x"04721013",
   565 => x"70842916",
   566 => x"51528812",
   567 => x"08802e89",
   568 => x"38fe5188",
   569 => x"12085271",
   570 => x"2d81fd51",
   571 => x"8bdd2db7",
   572 => x"a008812a",
   573 => x"70810651",
   574 => x"5271802e",
   575 => x"ad38b7fc",
   576 => x"08802e89",
   577 => x"38800bb7",
   578 => x"fc0c92aa",
   579 => x"04b7f808",
   580 => x"10b7f808",
   581 => x"05708429",
   582 => x"16515288",
   583 => x"1208802e",
   584 => x"8938fd51",
   585 => x"88120852",
   586 => x"712d81fa",
   587 => x"518bdd2d",
   588 => x"b7a00881",
   589 => x"2a708106",
   590 => x"51527180",
   591 => x"2eae38b7",
   592 => x"f808ff11",
   593 => x"5452b7fc",
   594 => x"08732588",
   595 => x"3872b7fc",
   596 => x"0c92ec04",
   597 => x"71101270",
   598 => x"84291651",
   599 => x"52881208",
   600 => x"802e8938",
   601 => x"fc518812",
   602 => x"0852712d",
   603 => x"b7fc0870",
   604 => x"53547380",
   605 => x"2e8a388c",
   606 => x"15ff1555",
   607 => x"5592f204",
   608 => x"820bb7b4",
   609 => x"0c718f06",
   610 => x"b7b00c81",
   611 => x"eb518bdd",
   612 => x"2db7a008",
   613 => x"812a7081",
   614 => x"06515271",
   615 => x"802ead38",
   616 => x"7408852e",
   617 => x"098106a4",
   618 => x"38881580",
   619 => x"f52dff05",
   620 => x"52718816",
   621 => x"81b72d71",
   622 => x"982b5271",
   623 => x"80258838",
   624 => x"800b8816",
   625 => x"81b72d74",
   626 => x"518e812d",
   627 => x"81f4518b",
   628 => x"dd2db7a0",
   629 => x"08812a70",
   630 => x"81065152",
   631 => x"71802eb3",
   632 => x"38740885",
   633 => x"2e098106",
   634 => x"aa388815",
   635 => x"80f52d81",
   636 => x"05527188",
   637 => x"1681b72d",
   638 => x"7181ff06",
   639 => x"8b1680f5",
   640 => x"2d545272",
   641 => x"72278738",
   642 => x"72881681",
   643 => x"b72d7451",
   644 => x"8e812d80",
   645 => x"da518bdd",
   646 => x"2db7a008",
   647 => x"812a7081",
   648 => x"06515271",
   649 => x"802e81a6",
   650 => x"38b7f408",
   651 => x"b7fc0855",
   652 => x"5373802e",
   653 => x"8a388c13",
   654 => x"ff155553",
   655 => x"94b10472",
   656 => x"08527182",
   657 => x"2ea63871",
   658 => x"82268938",
   659 => x"71812ea9",
   660 => x"3895ce04",
   661 => x"71832eb1",
   662 => x"3871842e",
   663 => x"09810680",
   664 => x"ed388813",
   665 => x"08518fcc",
   666 => x"2d95ce04",
   667 => x"b7fc0851",
   668 => x"88130852",
   669 => x"712d95ce",
   670 => x"04810b88",
   671 => x"14082bb5",
   672 => x"dc0832b5",
   673 => x"dc0c95a4",
   674 => x"04881380",
   675 => x"f52d8105",
   676 => x"8b1480f5",
   677 => x"2d535471",
   678 => x"74248338",
   679 => x"80547388",
   680 => x"1481b72d",
   681 => x"8eb12d95",
   682 => x"ce047508",
   683 => x"802ea238",
   684 => x"7508518b",
   685 => x"dd2db7a0",
   686 => x"08810652",
   687 => x"71802e8b",
   688 => x"38b7fc08",
   689 => x"51841608",
   690 => x"52712d88",
   691 => x"165675da",
   692 => x"38805480",
   693 => x"0bb7b40c",
   694 => x"738f06b7",
   695 => x"b00ca052",
   696 => x"73b7fc08",
   697 => x"2e098106",
   698 => x"9838b7f8",
   699 => x"08ff0574",
   700 => x"32700981",
   701 => x"05707207",
   702 => x"9f2a9171",
   703 => x"31515153",
   704 => x"53715182",
   705 => x"f92d8114",
   706 => x"548e7425",
   707 => x"c638b5e0",
   708 => x"085271b7",
   709 => x"a00c0298",
   710 => x"050d0402",
   711 => x"f4050dd4",
   712 => x"5281ff72",
   713 => x"0c710853",
   714 => x"81ff720c",
   715 => x"72882b83",
   716 => x"fe800672",
   717 => x"087081ff",
   718 => x"06515253",
   719 => x"81ff720c",
   720 => x"72710788",
   721 => x"2b720870",
   722 => x"81ff0651",
   723 => x"525381ff",
   724 => x"720c7271",
   725 => x"07882b72",
   726 => x"087081ff",
   727 => x"067207b7",
   728 => x"a00c5253",
   729 => x"028c050d",
   730 => x"0402f405",
   731 => x"0d747671",
   732 => x"81ff06d4",
   733 => x"0c5353b8",
   734 => x"84088538",
   735 => x"71892b52",
   736 => x"71982ad4",
   737 => x"0c71902a",
   738 => x"7081ff06",
   739 => x"d40c5171",
   740 => x"882a7081",
   741 => x"ff06d40c",
   742 => x"517181ff",
   743 => x"06d40c72",
   744 => x"902a7081",
   745 => x"ff06d40c",
   746 => x"51d40870",
   747 => x"81ff0651",
   748 => x"5182b8bf",
   749 => x"527081ff",
   750 => x"2e098106",
   751 => x"943881ff",
   752 => x"0bd40cd4",
   753 => x"087081ff",
   754 => x"06ff1454",
   755 => x"515171e5",
   756 => x"3870b7a0",
   757 => x"0c028c05",
   758 => x"0d0402fc",
   759 => x"050d81c7",
   760 => x"5181ff0b",
   761 => x"d40cff11",
   762 => x"51708025",
   763 => x"f4380284",
   764 => x"050d0402",
   765 => x"f4050d81",
   766 => x"ff0bd40c",
   767 => x"93538052",
   768 => x"87fc80c1",
   769 => x"5196e92d",
   770 => x"b7a0088b",
   771 => x"3881ff0b",
   772 => x"d40c8153",
   773 => x"98a00497",
   774 => x"da2dff13",
   775 => x"5372df38",
   776 => x"72b7a00c",
   777 => x"028c050d",
   778 => x"0402ec05",
   779 => x"0d810bb8",
   780 => x"840c8454",
   781 => x"d008708f",
   782 => x"2a708106",
   783 => x"51515372",
   784 => x"f33872d0",
   785 => x"0c97da2d",
   786 => x"b1fc5185",
   787 => x"fe2dd008",
   788 => x"708f2a70",
   789 => x"81065151",
   790 => x"5372f338",
   791 => x"810bd00c",
   792 => x"b1538052",
   793 => x"84d480c0",
   794 => x"5196e92d",
   795 => x"b7a00881",
   796 => x"2e933872",
   797 => x"822ebd38",
   798 => x"ff135372",
   799 => x"e538ff14",
   800 => x"5473ffb0",
   801 => x"3897da2d",
   802 => x"83aa5284",
   803 => x"9c80c851",
   804 => x"96e92db7",
   805 => x"a008812e",
   806 => x"09810692",
   807 => x"38969b2d",
   808 => x"b7a00883",
   809 => x"ffff0653",
   810 => x"7283aa2e",
   811 => x"9d3897f3",
   812 => x"2d99c504",
   813 => x"b2885185",
   814 => x"fe2d8053",
   815 => x"9b9304b2",
   816 => x"a05185fe",
   817 => x"2d80549a",
   818 => x"e50481ff",
   819 => x"0bd40cb1",
   820 => x"5497da2d",
   821 => x"8fcf5380",
   822 => x"5287fc80",
   823 => x"f75196e9",
   824 => x"2db7a008",
   825 => x"55b7a008",
   826 => x"812e0981",
   827 => x"069b3881",
   828 => x"ff0bd40c",
   829 => x"820a5284",
   830 => x"9c80e951",
   831 => x"96e92db7",
   832 => x"a008802e",
   833 => x"8d3897da",
   834 => x"2dff1353",
   835 => x"72c9389a",
   836 => x"d80481ff",
   837 => x"0bd40cb7",
   838 => x"a0085287",
   839 => x"fc80fa51",
   840 => x"96e92db7",
   841 => x"a008b138",
   842 => x"81ff0bd4",
   843 => x"0cd40853",
   844 => x"81ff0bd4",
   845 => x"0c81ff0b",
   846 => x"d40c81ff",
   847 => x"0bd40c81",
   848 => x"ff0bd40c",
   849 => x"72862a70",
   850 => x"81067656",
   851 => x"51537295",
   852 => x"38b7a008",
   853 => x"549ae504",
   854 => x"73822efe",
   855 => x"e238ff14",
   856 => x"5473feed",
   857 => x"3873b884",
   858 => x"0c738b38",
   859 => x"815287fc",
   860 => x"80d05196",
   861 => x"e92d81ff",
   862 => x"0bd40cd0",
   863 => x"08708f2a",
   864 => x"70810651",
   865 => x"515372f3",
   866 => x"3872d00c",
   867 => x"81ff0bd4",
   868 => x"0c815372",
   869 => x"b7a00c02",
   870 => x"94050d04",
   871 => x"02e8050d",
   872 => x"78558056",
   873 => x"81ff0bd4",
   874 => x"0cd00870",
   875 => x"8f2a7081",
   876 => x"06515153",
   877 => x"72f33882",
   878 => x"810bd00c",
   879 => x"81ff0bd4",
   880 => x"0c775287",
   881 => x"fc80d151",
   882 => x"96e92d80",
   883 => x"dbc6df54",
   884 => x"b7a00880",
   885 => x"2e8a38b2",
   886 => x"c05185fe",
   887 => x"2d9cb304",
   888 => x"81ff0bd4",
   889 => x"0cd40870",
   890 => x"81ff0651",
   891 => x"537281fe",
   892 => x"2e098106",
   893 => x"9d3880ff",
   894 => x"53969b2d",
   895 => x"b7a00875",
   896 => x"70840557",
   897 => x"0cff1353",
   898 => x"728025ed",
   899 => x"3881569c",
   900 => x"9804ff14",
   901 => x"5473c938",
   902 => x"81ff0bd4",
   903 => x"0c81ff0b",
   904 => x"d40cd008",
   905 => x"708f2a70",
   906 => x"81065151",
   907 => x"5372f338",
   908 => x"72d00c75",
   909 => x"b7a00c02",
   910 => x"98050d04",
   911 => x"02e8050d",
   912 => x"77797b58",
   913 => x"55558053",
   914 => x"727625a3",
   915 => x"38747081",
   916 => x"055680f5",
   917 => x"2d747081",
   918 => x"055680f5",
   919 => x"2d525271",
   920 => x"712e8638",
   921 => x"81519cf1",
   922 => x"04811353",
   923 => x"9cc80480",
   924 => x"5170b7a0",
   925 => x"0c029805",
   926 => x"0d0402ec",
   927 => x"050d7655",
   928 => x"74802ebb",
   929 => x"389a1580",
   930 => x"e02d51a9",
   931 => x"fa2db7a0",
   932 => x"08b7a008",
   933 => x"beb80cb7",
   934 => x"a0085454",
   935 => x"be940880",
   936 => x"2e993894",
   937 => x"1580e02d",
   938 => x"51a9fa2d",
   939 => x"b7a00890",
   940 => x"2b83fff0",
   941 => x"0a067075",
   942 => x"07515372",
   943 => x"beb80cbe",
   944 => x"b8085372",
   945 => x"802e9938",
   946 => x"be8c08fe",
   947 => x"147129be",
   948 => x"a00805be",
   949 => x"bc0c7084",
   950 => x"2bbe980c",
   951 => x"549e8604",
   952 => x"bea408be",
   953 => x"b80cbea8",
   954 => x"08bebc0c",
   955 => x"be940880",
   956 => x"2e8a38be",
   957 => x"8c08842b",
   958 => x"539e8204",
   959 => x"beac0884",
   960 => x"2b5372be",
   961 => x"980c0294",
   962 => x"050d0402",
   963 => x"d8050d80",
   964 => x"0bbe940c",
   965 => x"845498a9",
   966 => x"2db7a008",
   967 => x"802e9538",
   968 => x"b8885280",
   969 => x"519b9c2d",
   970 => x"b7a00880",
   971 => x"2e8638fe",
   972 => x"549ebc04",
   973 => x"ff145473",
   974 => x"8024db38",
   975 => x"738c38b2",
   976 => x"d05185fe",
   977 => x"2d7355a3",
   978 => x"c5048056",
   979 => x"810bbec0",
   980 => x"0c8853b2",
   981 => x"e452b8be",
   982 => x"519cbc2d",
   983 => x"b7a00876",
   984 => x"2e098106",
   985 => x"8738b7a0",
   986 => x"08bec00c",
   987 => x"8853b2f0",
   988 => x"52b8da51",
   989 => x"9cbc2db7",
   990 => x"a0088738",
   991 => x"b7a008be",
   992 => x"c00cbec0",
   993 => x"08802e80",
   994 => x"f638bbce",
   995 => x"0b80f52d",
   996 => x"bbcf0b80",
   997 => x"f52d7198",
   998 => x"2b71902b",
   999 => x"07bbd00b",
  1000 => x"80f52d70",
  1001 => x"882b7207",
  1002 => x"bbd10b80",
  1003 => x"f52d7107",
  1004 => x"bc860b80",
  1005 => x"f52dbc87",
  1006 => x"0b80f52d",
  1007 => x"71882b07",
  1008 => x"535f5452",
  1009 => x"5a565755",
  1010 => x"7381abaa",
  1011 => x"2e098106",
  1012 => x"8d387551",
  1013 => x"a9ca2db7",
  1014 => x"a008569f",
  1015 => x"eb047382",
  1016 => x"d4d52e87",
  1017 => x"38b2fc51",
  1018 => x"a0ac04b8",
  1019 => x"88527551",
  1020 => x"9b9c2db7",
  1021 => x"a00855b7",
  1022 => x"a008802e",
  1023 => x"83c73888",
  1024 => x"53b2f052",
  1025 => x"b8da519c",
  1026 => x"bc2db7a0",
  1027 => x"08893881",
  1028 => x"0bbe940c",
  1029 => x"a0b20488",
  1030 => x"53b2e452",
  1031 => x"b8be519c",
  1032 => x"bc2db7a0",
  1033 => x"08802e8a",
  1034 => x"38b39051",
  1035 => x"85fe2da1",
  1036 => x"8c04bc86",
  1037 => x"0b80f52d",
  1038 => x"547380d5",
  1039 => x"2e098106",
  1040 => x"80ca38bc",
  1041 => x"870b80f5",
  1042 => x"2d547381",
  1043 => x"aa2e0981",
  1044 => x"06ba3880",
  1045 => x"0bb8880b",
  1046 => x"80f52d56",
  1047 => x"547481e9",
  1048 => x"2e833881",
  1049 => x"547481eb",
  1050 => x"2e8c3880",
  1051 => x"5573752e",
  1052 => x"09810682",
  1053 => x"d038b893",
  1054 => x"0b80f52d",
  1055 => x"55748d38",
  1056 => x"b8940b80",
  1057 => x"f52d5473",
  1058 => x"822e8638",
  1059 => x"8055a3c5",
  1060 => x"04b8950b",
  1061 => x"80f52d70",
  1062 => x"be8c0cff",
  1063 => x"05be900c",
  1064 => x"b8960b80",
  1065 => x"f52db897",
  1066 => x"0b80f52d",
  1067 => x"58760577",
  1068 => x"82802905",
  1069 => x"70be9c0c",
  1070 => x"b8980b80",
  1071 => x"f52d70be",
  1072 => x"b00cbe94",
  1073 => x"08595758",
  1074 => x"76802e81",
  1075 => x"a3388853",
  1076 => x"b2f052b8",
  1077 => x"da519cbc",
  1078 => x"2db7a008",
  1079 => x"81e738be",
  1080 => x"8c087084",
  1081 => x"2bbe980c",
  1082 => x"70beac0c",
  1083 => x"b8ad0b80",
  1084 => x"f52db8ac",
  1085 => x"0b80f52d",
  1086 => x"71828029",
  1087 => x"05b8ae0b",
  1088 => x"80f52d70",
  1089 => x"84808029",
  1090 => x"12b8af0b",
  1091 => x"80f52d70",
  1092 => x"81800a29",
  1093 => x"1270beb4",
  1094 => x"0cbeb008",
  1095 => x"7129be9c",
  1096 => x"080570be",
  1097 => x"a00cb8b5",
  1098 => x"0b80f52d",
  1099 => x"b8b40b80",
  1100 => x"f52d7182",
  1101 => x"802905b8",
  1102 => x"b60b80f5",
  1103 => x"2d708480",
  1104 => x"802912b8",
  1105 => x"b70b80f5",
  1106 => x"2d70982b",
  1107 => x"81f00a06",
  1108 => x"720570be",
  1109 => x"a40cfe11",
  1110 => x"7e297705",
  1111 => x"bea80c52",
  1112 => x"59524354",
  1113 => x"5e515259",
  1114 => x"525d5759",
  1115 => x"57a3be04",
  1116 => x"b89a0b80",
  1117 => x"f52db899",
  1118 => x"0b80f52d",
  1119 => x"71828029",
  1120 => x"0570be98",
  1121 => x"0c70a029",
  1122 => x"83ff0570",
  1123 => x"892a70be",
  1124 => x"ac0cb89f",
  1125 => x"0b80f52d",
  1126 => x"b89e0b80",
  1127 => x"f52d7182",
  1128 => x"80290570",
  1129 => x"beb40c7b",
  1130 => x"71291e70",
  1131 => x"bea80c7d",
  1132 => x"bea40c73",
  1133 => x"05bea00c",
  1134 => x"555e5151",
  1135 => x"55558051",
  1136 => x"9cfa2d81",
  1137 => x"5574b7a0",
  1138 => x"0c02a805",
  1139 => x"0d0402ec",
  1140 => x"050d7670",
  1141 => x"872c7180",
  1142 => x"ff065556",
  1143 => x"54be9408",
  1144 => x"8a387388",
  1145 => x"2c7481ff",
  1146 => x"065455b8",
  1147 => x"8852be9c",
  1148 => x"0815519b",
  1149 => x"9c2db7a0",
  1150 => x"0854b7a0",
  1151 => x"08802eb3",
  1152 => x"38be9408",
  1153 => x"802e9838",
  1154 => x"728429b8",
  1155 => x"88057008",
  1156 => x"5253a9ca",
  1157 => x"2db7a008",
  1158 => x"f00a0653",
  1159 => x"a4b10472",
  1160 => x"10b88805",
  1161 => x"7080e02d",
  1162 => x"5253a9fa",
  1163 => x"2db7a008",
  1164 => x"53725473",
  1165 => x"b7a00c02",
  1166 => x"94050d04",
  1167 => x"02e0050d",
  1168 => x"7970842c",
  1169 => x"bebc0805",
  1170 => x"718f0652",
  1171 => x"55537289",
  1172 => x"38b88852",
  1173 => x"73519b9c",
  1174 => x"2d72a029",
  1175 => x"b8880554",
  1176 => x"807480f5",
  1177 => x"2d565374",
  1178 => x"732e8338",
  1179 => x"81537481",
  1180 => x"e52e81ef",
  1181 => x"38817074",
  1182 => x"06545872",
  1183 => x"802e81e3",
  1184 => x"388b1480",
  1185 => x"f52d7083",
  1186 => x"2a790658",
  1187 => x"56769838",
  1188 => x"b5e40853",
  1189 => x"72883872",
  1190 => x"bc880b81",
  1191 => x"b72d76b5",
  1192 => x"e40c7353",
  1193 => x"a6e50475",
  1194 => x"8f2e0981",
  1195 => x"0681b438",
  1196 => x"749f068d",
  1197 => x"29bbfb11",
  1198 => x"51538114",
  1199 => x"80f52d73",
  1200 => x"70810555",
  1201 => x"81b72d83",
  1202 => x"1480f52d",
  1203 => x"73708105",
  1204 => x"5581b72d",
  1205 => x"851480f5",
  1206 => x"2d737081",
  1207 => x"055581b7",
  1208 => x"2d871480",
  1209 => x"f52d7370",
  1210 => x"81055581",
  1211 => x"b72d8914",
  1212 => x"80f52d73",
  1213 => x"70810555",
  1214 => x"81b72d8e",
  1215 => x"1480f52d",
  1216 => x"73708105",
  1217 => x"5581b72d",
  1218 => x"901480f5",
  1219 => x"2d737081",
  1220 => x"055581b7",
  1221 => x"2d921480",
  1222 => x"f52d7370",
  1223 => x"81055581",
  1224 => x"b72d9414",
  1225 => x"80f52d73",
  1226 => x"70810555",
  1227 => x"81b72d96",
  1228 => x"1480f52d",
  1229 => x"73708105",
  1230 => x"5581b72d",
  1231 => x"981480f5",
  1232 => x"2d737081",
  1233 => x"055581b7",
  1234 => x"2d9c1480",
  1235 => x"f52d7370",
  1236 => x"81055581",
  1237 => x"b72d9e14",
  1238 => x"80f52d73",
  1239 => x"81b72d77",
  1240 => x"b5e40c80",
  1241 => x"5372b7a0",
  1242 => x"0c02a005",
  1243 => x"0d0402cc",
  1244 => x"050d7e60",
  1245 => x"5e5a800b",
  1246 => x"beb808be",
  1247 => x"bc08595c",
  1248 => x"568058be",
  1249 => x"9808782e",
  1250 => x"81ae3877",
  1251 => x"8f06a017",
  1252 => x"5754738f",
  1253 => x"38b88852",
  1254 => x"76518117",
  1255 => x"579b9c2d",
  1256 => x"b8885680",
  1257 => x"7680f52d",
  1258 => x"56547474",
  1259 => x"2e833881",
  1260 => x"547481e5",
  1261 => x"2e80f638",
  1262 => x"81707506",
  1263 => x"555c7380",
  1264 => x"2e80ea38",
  1265 => x"8b1680f5",
  1266 => x"2d980659",
  1267 => x"7880de38",
  1268 => x"8b537c52",
  1269 => x"75519cbc",
  1270 => x"2db7a008",
  1271 => x"80cf389c",
  1272 => x"160851a9",
  1273 => x"ca2db7a0",
  1274 => x"08841b0c",
  1275 => x"9a1680e0",
  1276 => x"2d51a9fa",
  1277 => x"2db7a008",
  1278 => x"b7a00888",
  1279 => x"1c0cb7a0",
  1280 => x"085555be",
  1281 => x"9408802e",
  1282 => x"98389416",
  1283 => x"80e02d51",
  1284 => x"a9fa2db7",
  1285 => x"a008902b",
  1286 => x"83fff00a",
  1287 => x"06701651",
  1288 => x"5473881b",
  1289 => x"0c787a0c",
  1290 => x"7b54a8ee",
  1291 => x"04811858",
  1292 => x"be980878",
  1293 => x"26fed438",
  1294 => x"be940880",
  1295 => x"2eae387a",
  1296 => x"51a3ce2d",
  1297 => x"b7a008b7",
  1298 => x"a00880ff",
  1299 => x"fffff806",
  1300 => x"555b7380",
  1301 => x"fffffff8",
  1302 => x"2e9238b7",
  1303 => x"a008fe05",
  1304 => x"be8c0829",
  1305 => x"bea00805",
  1306 => x"57a78104",
  1307 => x"805473b7",
  1308 => x"a00c02b4",
  1309 => x"050d0402",
  1310 => x"f4050d74",
  1311 => x"70088105",
  1312 => x"710c7008",
  1313 => x"be900806",
  1314 => x"5353718e",
  1315 => x"38881308",
  1316 => x"51a3ce2d",
  1317 => x"b7a00888",
  1318 => x"140c810b",
  1319 => x"b7a00c02",
  1320 => x"8c050d04",
  1321 => x"02f0050d",
  1322 => x"75881108",
  1323 => x"fe05be8c",
  1324 => x"0829bea0",
  1325 => x"08117208",
  1326 => x"be900806",
  1327 => x"05795553",
  1328 => x"54549b9c",
  1329 => x"2d029005",
  1330 => x"0d0402f4",
  1331 => x"050d7470",
  1332 => x"882a83fe",
  1333 => x"80067072",
  1334 => x"982a0772",
  1335 => x"882b87fc",
  1336 => x"80800673",
  1337 => x"982b81f0",
  1338 => x"0a067173",
  1339 => x"0707b7a0",
  1340 => x"0c565153",
  1341 => x"51028c05",
  1342 => x"0d0402f8",
  1343 => x"050d028e",
  1344 => x"0580f52d",
  1345 => x"74882b07",
  1346 => x"7083ffff",
  1347 => x"06b7a00c",
  1348 => x"51028805",
  1349 => x"0d0402f4",
  1350 => x"050d7476",
  1351 => x"78535452",
  1352 => x"80712597",
  1353 => x"38727081",
  1354 => x"055480f5",
  1355 => x"2d727081",
  1356 => x"055481b7",
  1357 => x"2dff1151",
  1358 => x"70eb3880",
  1359 => x"7281b72d",
  1360 => x"028c050d",
  1361 => x"0402e805",
  1362 => x"0d775680",
  1363 => x"70565473",
  1364 => x"7624b138",
  1365 => x"be980874",
  1366 => x"2eaa3873",
  1367 => x"51a4bc2d",
  1368 => x"b7a008b7",
  1369 => x"a0080981",
  1370 => x"0570b7a0",
  1371 => x"08079f2a",
  1372 => x"77058117",
  1373 => x"57575353",
  1374 => x"74762488",
  1375 => x"38be9808",
  1376 => x"7426d838",
  1377 => x"72b7a00c",
  1378 => x"0298050d",
  1379 => x"0402f005",
  1380 => x"0db79c08",
  1381 => x"1651aac5",
  1382 => x"2db7a008",
  1383 => x"802e9b38",
  1384 => x"8b53b7a0",
  1385 => x"0852bc88",
  1386 => x"51aa962d",
  1387 => x"bec40854",
  1388 => x"73802e86",
  1389 => x"38bc8851",
  1390 => x"732d0290",
  1391 => x"050d0402",
  1392 => x"dc050d80",
  1393 => x"705a5574",
  1394 => x"b79c0825",
  1395 => x"af38be98",
  1396 => x"08752ea8",
  1397 => x"387851a4",
  1398 => x"bc2db7a0",
  1399 => x"08098105",
  1400 => x"70b7a008",
  1401 => x"079f2a76",
  1402 => x"05811b5b",
  1403 => x"565474b7",
  1404 => x"9c082588",
  1405 => x"38be9808",
  1406 => x"7926da38",
  1407 => x"805578be",
  1408 => x"98082781",
  1409 => x"cd387851",
  1410 => x"a4bc2db7",
  1411 => x"a008802e",
  1412 => x"81a238b7",
  1413 => x"a0088b05",
  1414 => x"80f52d70",
  1415 => x"842a7081",
  1416 => x"06771078",
  1417 => x"842bbc88",
  1418 => x"0b80f52d",
  1419 => x"5c5c5351",
  1420 => x"55567380",
  1421 => x"2e80c638",
  1422 => x"7416822b",
  1423 => x"adf50bb5",
  1424 => x"f0120c54",
  1425 => x"77753110",
  1426 => x"bec81155",
  1427 => x"56907470",
  1428 => x"81055681",
  1429 => x"b72da074",
  1430 => x"81b72d76",
  1431 => x"81ff0681",
  1432 => x"16585473",
  1433 => x"802e8938",
  1434 => x"9c53bc88",
  1435 => x"52acf604",
  1436 => x"8b53b7a0",
  1437 => x"0852beca",
  1438 => x"1651adac",
  1439 => x"04741682",
  1440 => x"2bab8d0b",
  1441 => x"b5f0120c",
  1442 => x"547681ff",
  1443 => x"06811658",
  1444 => x"5473802e",
  1445 => x"89389c53",
  1446 => x"bc8852ad",
  1447 => x"a4048b53",
  1448 => x"b7a00852",
  1449 => x"77753110",
  1450 => x"bec80551",
  1451 => x"7655aa96",
  1452 => x"2dadc704",
  1453 => x"74902975",
  1454 => x"317010be",
  1455 => x"c8055154",
  1456 => x"b7a00874",
  1457 => x"81b72d81",
  1458 => x"1959748b",
  1459 => x"24a238ab",
  1460 => x"fe047490",
  1461 => x"29753170",
  1462 => x"10bec805",
  1463 => x"8c773157",
  1464 => x"51548074",
  1465 => x"81b72d9e",
  1466 => x"14ff1656",
  1467 => x"5474f338",
  1468 => x"02a4050d",
  1469 => x"0402fc05",
  1470 => x"0db79c08",
  1471 => x"1351aac5",
  1472 => x"2db7a008",
  1473 => x"802e8838",
  1474 => x"b7a00851",
  1475 => x"9cfa2d80",
  1476 => x"0bb79c0c",
  1477 => x"abbf2d8e",
  1478 => x"b12d0284",
  1479 => x"050d0402",
  1480 => x"fc050d72",
  1481 => x"5170fd2e",
  1482 => x"ad3870fd",
  1483 => x"248a3870",
  1484 => x"fc2e80c4",
  1485 => x"38af8004",
  1486 => x"70fe2eb1",
  1487 => x"3870ff2e",
  1488 => x"098106bc",
  1489 => x"38b79c08",
  1490 => x"5170802e",
  1491 => x"b338ff11",
  1492 => x"b79c0caf",
  1493 => x"8004b79c",
  1494 => x"08f00570",
  1495 => x"b79c0c51",
  1496 => x"7080259c",
  1497 => x"38800bb7",
  1498 => x"9c0caf80",
  1499 => x"04b79c08",
  1500 => x"8105b79c",
  1501 => x"0caf8004",
  1502 => x"b79c0890",
  1503 => x"05b79c0c",
  1504 => x"abbf2d8e",
  1505 => x"b12d0284",
  1506 => x"050d0402",
  1507 => x"fc050d80",
  1508 => x"0bb79c0c",
  1509 => x"abbf2d8d",
  1510 => x"c82db7a0",
  1511 => x"08b78c0c",
  1512 => x"b5e8518f",
  1513 => x"cc2d0284",
  1514 => x"050d0471",
  1515 => x"bec40c04",
  1516 => x"00ffffff",
  1517 => x"ff00ffff",
  1518 => x"ffff00ff",
  1519 => x"ffffff00",
  1520 => x"2020203d",
  1521 => x"52616d70",
  1522 => x"61205669",
  1523 => x"64656f70",
  1524 => x"61633d20",
  1525 => x"20202000",
  1526 => x"20202020",
  1527 => x"20202020",
  1528 => x"20202020",
  1529 => x"20202020",
  1530 => x"20202020",
  1531 => x"20202000",
  1532 => x"52657365",
  1533 => x"74000000",
  1534 => x"43617267",
  1535 => x"61722043",
  1536 => x"61727475",
  1537 => x"63686f2f",
  1538 => x"466f6e74",
  1539 => x"20100000",
  1540 => x"45786974",
  1541 => x"00000000",
  1542 => x"54562043",
  1543 => x"6f6c6f72",
  1544 => x"00000000",
  1545 => x"54562042",
  1546 => x"2f570000",
  1547 => x"4f647973",
  1548 => x"73657932",
  1549 => x"00000000",
  1550 => x"56696465",
  1551 => x"6f706163",
  1552 => x"00000000",
  1553 => x"436f6d70",
  1554 => x"6f736974",
  1555 => x"65000000",
  1556 => x"52474200",
  1557 => x"54686520",
  1558 => x"566f6963",
  1559 => x"65204f66",
  1560 => x"66000000",
  1561 => x"54686520",
  1562 => x"566f6963",
  1563 => x"65204f6e",
  1564 => x"00000000",
  1565 => x"53776170",
  1566 => x"204a6f79",
  1567 => x"204f6666",
  1568 => x"00000000",
  1569 => x"53776170",
  1570 => x"206a6f79",
  1571 => x"204f6e00",
  1572 => x"5363616e",
  1573 => x"6c696e65",
  1574 => x"73204e6f",
  1575 => x"6e650000",
  1576 => x"5363616e",
  1577 => x"6c696e65",
  1578 => x"73204352",
  1579 => x"54203235",
  1580 => x"25000000",
  1581 => x"5363616e",
  1582 => x"6c696e65",
  1583 => x"73204352",
  1584 => x"54203530",
  1585 => x"25000000",
  1586 => x"5363616e",
  1587 => x"6c696e65",
  1588 => x"73204352",
  1589 => x"54203735",
  1590 => x"25000000",
  1591 => x"43617267",
  1592 => x"61204661",
  1593 => x"6c6c6964",
  1594 => x"61000000",
  1595 => x"4f4b0000",
  1596 => x"16200000",
  1597 => x"14200000",
  1598 => x"15200000",
  1599 => x"53442069",
  1600 => x"6e69742e",
  1601 => x"2e2e0a00",
  1602 => x"53442063",
  1603 => x"61726420",
  1604 => x"72657365",
  1605 => x"74206661",
  1606 => x"696c6564",
  1607 => x"210a0000",
  1608 => x"53444843",
  1609 => x"20657272",
  1610 => x"6f72210a",
  1611 => x"00000000",
  1612 => x"57726974",
  1613 => x"65206661",
  1614 => x"696c6564",
  1615 => x"0a000000",
  1616 => x"52656164",
  1617 => x"20666169",
  1618 => x"6c65640a",
  1619 => x"00000000",
  1620 => x"43617264",
  1621 => x"20696e69",
  1622 => x"74206661",
  1623 => x"696c6564",
  1624 => x"0a000000",
  1625 => x"46415431",
  1626 => x"36202020",
  1627 => x"00000000",
  1628 => x"46415433",
  1629 => x"32202020",
  1630 => x"00000000",
  1631 => x"4e6f2070",
  1632 => x"61727469",
  1633 => x"74696f6e",
  1634 => x"20736967",
  1635 => x"0a000000",
  1636 => x"42616420",
  1637 => x"70617274",
  1638 => x"0a000000",
  1639 => x"4261636b",
  1640 => x"00000000",
  1641 => x"00000002",
  1642 => x"00000002",
  1643 => x"000017c0",
  1644 => x"00000000",
  1645 => x"00000002",
  1646 => x"000017d8",
  1647 => x"00000000",
  1648 => x"00000002",
  1649 => x"000017f0",
  1650 => x"0000034e",
  1651 => x"00000003",
  1652 => x"00001a60",
  1653 => x"00000004",
  1654 => x"00000003",
  1655 => x"00001a58",
  1656 => x"00000002",
  1657 => x"00000003",
  1658 => x"00001a50",
  1659 => x"00000002",
  1660 => x"00000003",
  1661 => x"00001a48",
  1662 => x"00000002",
  1663 => x"00000003",
  1664 => x"00001a40",
  1665 => x"00000002",
  1666 => x"00000003",
  1667 => x"00001a38",
  1668 => x"00000002",
  1669 => x"00000002",
  1670 => x"000017f8",
  1671 => x"0000178b",
  1672 => x"00000002",
  1673 => x"00001810",
  1674 => x"000006cf",
  1675 => x"00000000",
  1676 => x"00000000",
  1677 => x"00000000",
  1678 => x"00001818",
  1679 => x"00001824",
  1680 => x"0000182c",
  1681 => x"00001838",
  1682 => x"00001844",
  1683 => x"00001850",
  1684 => x"00001854",
  1685 => x"00001864",
  1686 => x"00001874",
  1687 => x"00001884",
  1688 => x"00001890",
  1689 => x"000018a0",
  1690 => x"000018b4",
  1691 => x"000018c8",
  1692 => x"00000004",
  1693 => x"000018dc",
  1694 => x"00001a70",
  1695 => x"00000004",
  1696 => x"000018ec",
  1697 => x"000019a8",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000000",
  1708 => x"00000000",
  1709 => x"00000000",
  1710 => x"00000000",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"00000000",
  1715 => x"00000000",
  1716 => x"00000000",
  1717 => x"00000000",
  1718 => x"00000000",
  1719 => x"00000000",
  1720 => x"00000000",
  1721 => x"00000000",
  1722 => x"00000002",
  1723 => x"00001f48",
  1724 => x"0000158d",
  1725 => x"00000002",
  1726 => x"00001f66",
  1727 => x"0000158d",
  1728 => x"00000002",
  1729 => x"00001f84",
  1730 => x"0000158d",
  1731 => x"00000002",
  1732 => x"00001fa2",
  1733 => x"0000158d",
  1734 => x"00000002",
  1735 => x"00001fc0",
  1736 => x"0000158d",
  1737 => x"00000002",
  1738 => x"00001fde",
  1739 => x"0000158d",
  1740 => x"00000002",
  1741 => x"00001ffc",
  1742 => x"0000158d",
  1743 => x"00000002",
  1744 => x"0000201a",
  1745 => x"0000158d",
  1746 => x"00000002",
  1747 => x"00002038",
  1748 => x"0000158d",
  1749 => x"00000002",
  1750 => x"00002056",
  1751 => x"0000158d",
  1752 => x"00000002",
  1753 => x"00002074",
  1754 => x"0000158d",
  1755 => x"00000002",
  1756 => x"00002092",
  1757 => x"0000158d",
  1758 => x"00000002",
  1759 => x"000020b0",
  1760 => x"0000158d",
  1761 => x"00000004",
  1762 => x"0000199c",
  1763 => x"00000000",
  1764 => x"00000000",
  1765 => x"00000000",
  1766 => x"0000171f",
  1767 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

