-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b80d1",
     9 => x"c0080b0b",
    10 => x"80d1c408",
    11 => x"0b0b80d1",
    12 => x"c8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b80",
    15 => x"d1c80c0b",
    16 => x"0b80d1c4",
    17 => x"0c0b0b80",
    18 => x"d1c00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bbdbc",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"80d1c070",
    57 => x"80dbfc27",
    58 => x"8b388071",
    59 => x"70840553",
    60 => x"0c81e304",
    61 => x"8c518aa2",
    62 => x"0402fc05",
    63 => x"0df88051",
    64 => x"8f0b80d1",
    65 => x"d00c9f0b",
    66 => x"80d1d40c",
    67 => x"a0717081",
    68 => x"05533480",
    69 => x"d1d408ff",
    70 => x"0580d1d4",
    71 => x"0c80d1d4",
    72 => x"088025e8",
    73 => x"3880d1d0",
    74 => x"08ff0580",
    75 => x"d1d00c80",
    76 => x"d1d00880",
    77 => x"25d03880",
    78 => x"0b80d1d4",
    79 => x"0c800b80",
    80 => x"d1d00c02",
    81 => x"84050d04",
    82 => x"02f0050d",
    83 => x"f88053f8",
    84 => x"a05483bf",
    85 => x"52737081",
    86 => x"05553351",
    87 => x"70737081",
    88 => x"055534ff",
    89 => x"12527180",
    90 => x"25eb38fb",
    91 => x"c0539f52",
    92 => x"a0737081",
    93 => x"055534ff",
    94 => x"12527180",
    95 => x"25f23802",
    96 => x"90050d04",
    97 => x"02f4050d",
    98 => x"74538e0b",
    99 => x"80d1d008",
   100 => x"25913882",
   101 => x"c82d80d1",
   102 => x"d008ff05",
   103 => x"80d1d00c",
   104 => x"838a0480",
   105 => x"d1d00880",
   106 => x"d1d40853",
   107 => x"51728a2e",
   108 => x"098106be",
   109 => x"38715171",
   110 => x"9f24a438",
   111 => x"80d1d008",
   112 => x"a02911f8",
   113 => x"80115151",
   114 => x"a0713480",
   115 => x"d1d40881",
   116 => x"0580d1d4",
   117 => x"0c80d1d4",
   118 => x"08519f71",
   119 => x"25de3880",
   120 => x"0b80d1d4",
   121 => x"0c80d1d0",
   122 => x"08810580",
   123 => x"d1d00c84",
   124 => x"880470a0",
   125 => x"2912f880",
   126 => x"11515172",
   127 => x"713480d1",
   128 => x"d4088105",
   129 => x"80d1d40c",
   130 => x"80d1d408",
   131 => x"a02e0981",
   132 => x"06913880",
   133 => x"0b80d1d4",
   134 => x"0c80d1d0",
   135 => x"08810580",
   136 => x"d1d00c02",
   137 => x"8c050d04",
   138 => x"02e8050d",
   139 => x"77795656",
   140 => x"880bfc16",
   141 => x"77712c8f",
   142 => x"06545254",
   143 => x"80537272",
   144 => x"25953871",
   145 => x"53fbe014",
   146 => x"51877134",
   147 => x"8114ff14",
   148 => x"545472f1",
   149 => x"387153f9",
   150 => x"1576712c",
   151 => x"87065351",
   152 => x"71802e8b",
   153 => x"38fbe014",
   154 => x"51717134",
   155 => x"81145472",
   156 => x"8e249538",
   157 => x"8f733153",
   158 => x"fbe01451",
   159 => x"a0713481",
   160 => x"14ff1454",
   161 => x"5472f138",
   162 => x"0298050d",
   163 => x"0402ec05",
   164 => x"0d800b80",
   165 => x"d1d80cf6",
   166 => x"8c08f690",
   167 => x"0871882c",
   168 => x"565381ff",
   169 => x"06537373",
   170 => x"25893872",
   171 => x"54820b80",
   172 => x"d1d80c71",
   173 => x"882c7281",
   174 => x"ff065355",
   175 => x"7472258d",
   176 => x"387180d1",
   177 => x"d8088407",
   178 => x"80d1d80c",
   179 => x"5573842b",
   180 => x"75832b56",
   181 => x"5485bc74",
   182 => x"258f3882",
   183 => x"0b0b0b80",
   184 => x"c8f80c80",
   185 => x"d05385f3",
   186 => x"04810b0b",
   187 => x"0b80c8f8",
   188 => x"0cbc530b",
   189 => x"0b80c8f8",
   190 => x"0881712b",
   191 => x"ff05f688",
   192 => x"0cfc0875",
   193 => x"7531ffb0",
   194 => x"05ff1371",
   195 => x"712cff94",
   196 => x"1a709f2a",
   197 => x"1170812c",
   198 => x"80d1d808",
   199 => x"52545153",
   200 => x"57535152",
   201 => x"5276802e",
   202 => x"85387081",
   203 => x"075170f6",
   204 => x"940c7209",
   205 => x"8105f680",
   206 => x"0c710981",
   207 => x"05f6840c",
   208 => x"0294050d",
   209 => x"0402f405",
   210 => x"0d745372",
   211 => x"70810554",
   212 => x"80f52d52",
   213 => x"71802e89",
   214 => x"38715183",
   215 => x"842d86cb",
   216 => x"04810b80",
   217 => x"d1c00c02",
   218 => x"8c050d04",
   219 => x"02fc050d",
   220 => x"81808051",
   221 => x"c0115170",
   222 => x"fb380284",
   223 => x"050d0402",
   224 => x"fc050dec",
   225 => x"5183710c",
   226 => x"86ec2d82",
   227 => x"710c0284",
   228 => x"050d0402",
   229 => x"fc050d84",
   230 => x"bf5186ec",
   231 => x"2dff1151",
   232 => x"708025f6",
   233 => x"38028405",
   234 => x"0d040402",
   235 => x"fc050d92",
   236 => x"c92d80d1",
   237 => x"c00880ce",
   238 => x"fc0c80cd",
   239 => x"d8519581",
   240 => x"2d028405",
   241 => x"0d0402fc",
   242 => x"050d92c9",
   243 => x"2d80d1c0",
   244 => x"0880cdc8",
   245 => x"0c80cca4",
   246 => x"5195812d",
   247 => x"0284050d",
   248 => x"0402dc05",
   249 => x"0d7a5580",
   250 => x"59840bec",
   251 => x"0c80c980",
   252 => x"085380c8",
   253 => x"fc08812e",
   254 => x"0981068c",
   255 => x"38728280",
   256 => x"0780c980",
   257 => x"0c889304",
   258 => x"72828007",
   259 => x"82803280",
   260 => x"c9800c80",
   261 => x"c98008fc",
   262 => x"0c86ec2d",
   263 => x"745280d1",
   264 => x"dc51b3f8",
   265 => x"2d80d1c0",
   266 => x"08802e81",
   267 => x"ae3880d1",
   268 => x"e0085480",
   269 => x"5673852e",
   270 => x"098106a5",
   271 => x"38745186",
   272 => x"c52d8793",
   273 => x"2d87932d",
   274 => x"87932d87",
   275 => x"932d8793",
   276 => x"2d87932d",
   277 => x"80d1e808",
   278 => x"5195812d",
   279 => x"81538a98",
   280 => x"0473f80c",
   281 => x"a50bec0c",
   282 => x"87932d84",
   283 => x"0bec0c75",
   284 => x"ff155758",
   285 => x"75802e8b",
   286 => x"38811876",
   287 => x"812a5758",
   288 => x"88f404f7",
   289 => x"18588159",
   290 => x"80742580",
   291 => x"ce387752",
   292 => x"755184a8",
   293 => x"2d80d2b4",
   294 => x"5280d1dc",
   295 => x"51b6c52d",
   296 => x"80d1c008",
   297 => x"802e9b38",
   298 => x"80d2b457",
   299 => x"83fc5576",
   300 => x"70840558",
   301 => x"08e80cfc",
   302 => x"15557480",
   303 => x"25f13889",
   304 => x"ca0480d1",
   305 => x"c0085984",
   306 => x"805480d1",
   307 => x"dc51b695",
   308 => x"2dfc8014",
   309 => x"81175754",
   310 => x"89880480",
   311 => x"c8fc0853",
   312 => x"72893872",
   313 => x"5186ff2d",
   314 => x"8a820480",
   315 => x"0b80c8fc",
   316 => x"0c80c980",
   317 => x"08828007",
   318 => x"82803270",
   319 => x"80c9800c",
   320 => x"fc0c7880",
   321 => x"2e893880",
   322 => x"d1e80851",
   323 => x"8a930480",
   324 => x"cc805195",
   325 => x"812d7853",
   326 => x"7280d1c0",
   327 => x"0c02a405",
   328 => x"0d0402e4",
   329 => x"050d900b",
   330 => x"80c9800c",
   331 => x"805186ff",
   332 => x"2d840bec",
   333 => x"0c92992d",
   334 => x"8ec42d81",
   335 => x"f92d8353",
   336 => x"91fc2d81",
   337 => x"51858d2d",
   338 => x"ff135372",
   339 => x"8025f138",
   340 => x"840bec0c",
   341 => x"80c7ac51",
   342 => x"86c52daa",
   343 => x"b02d80d1",
   344 => x"c008802e",
   345 => x"83c73881",
   346 => x"0bec0c84",
   347 => x"0bec0cbd",
   348 => x"cc5280d1",
   349 => x"dc51b3f8",
   350 => x"2d80d1c0",
   351 => x"08802e80",
   352 => x"cb3880d2",
   353 => x"b45280d1",
   354 => x"dc51b6c5",
   355 => x"2d80d1c0",
   356 => x"08802eb8",
   357 => x"3880d2b4",
   358 => x"0b80f52d",
   359 => x"80cfec0c",
   360 => x"80d2b50b",
   361 => x"80f52d80",
   362 => x"cff00c80",
   363 => x"d2b60b80",
   364 => x"f52d80cf",
   365 => x"f40c80d2",
   366 => x"b70b80f5",
   367 => x"2d80cff8",
   368 => x"0c80d2b8",
   369 => x"0b80f52d",
   370 => x"80cffc0c",
   371 => x"bddc5280",
   372 => x"d1dc51b3",
   373 => x"f82d80d1",
   374 => x"c008802e",
   375 => x"80cb3880",
   376 => x"d2b45280",
   377 => x"d1dc51b6",
   378 => x"c52d80d1",
   379 => x"c008802e",
   380 => x"b83880d2",
   381 => x"b40b80f5",
   382 => x"2d80cfd8",
   383 => x"0c80d2b5",
   384 => x"0b80f52d",
   385 => x"80cfdc0c",
   386 => x"80d2b60b",
   387 => x"80f52d80",
   388 => x"cfe00c80",
   389 => x"d2b70b80",
   390 => x"f52d80cf",
   391 => x"e40c80d2",
   392 => x"b80b80f5",
   393 => x"2d80cfe8",
   394 => x"0c87e151",
   395 => x"bdb52d80",
   396 => x"c9800880",
   397 => x"cfd40c80",
   398 => x"c98008fc",
   399 => x"0c80d294",
   400 => x"08882a70",
   401 => x"81065153",
   402 => x"72802e8c",
   403 => x"3880cacc",
   404 => x"0b80d1e8",
   405 => x"0c8ce004",
   406 => x"80c9840b",
   407 => x"80d1e80c",
   408 => x"80d1e808",
   409 => x"5195812d",
   410 => x"860b80d2",
   411 => x"a80c92d2",
   412 => x"2d8ed02d",
   413 => x"95942d80",
   414 => x"d1c00880",
   415 => x"d1e80880",
   416 => x"e81180f5",
   417 => x"2d70842b",
   418 => x"7080c980",
   419 => x"0c80f413",
   420 => x"80f52d70",
   421 => x"852b7207",
   422 => x"7080c980",
   423 => x"0c80d294",
   424 => x"08882a70",
   425 => x"81068180",
   426 => x"1780f52d",
   427 => x"80cfd408",
   428 => x"55575153",
   429 => x"535a5657",
   430 => x"55577280",
   431 => x"2e8b3873",
   432 => x"822b87fc",
   433 => x"06538dd1",
   434 => x"0473892b",
   435 => x"87fc8006",
   436 => x"53747307",
   437 => x"80c9800c",
   438 => x"75810653",
   439 => x"72802e8b",
   440 => x"3880c980",
   441 => x"08810780",
   442 => x"c9800c75",
   443 => x"812a7081",
   444 => x"06515372",
   445 => x"802e8b38",
   446 => x"80c98008",
   447 => x"820780c9",
   448 => x"800c7582",
   449 => x"2a708106",
   450 => x"51537280",
   451 => x"2e8c3880",
   452 => x"c9800881",
   453 => x"800780c9",
   454 => x"800c80c9",
   455 => x"8008fc0c",
   456 => x"86537683",
   457 => x"38845372",
   458 => x"ec0c8cf1",
   459 => x"04800b80",
   460 => x"d1c00c02",
   461 => x"9c050d04",
   462 => x"71980c04",
   463 => x"ffb00880",
   464 => x"d1c00c04",
   465 => x"810bffb0",
   466 => x"0c04800b",
   467 => x"ffb00c04",
   468 => x"02f4050d",
   469 => x"8fde0480",
   470 => x"d1c00881",
   471 => x"f02e0981",
   472 => x"068a3881",
   473 => x"0b80cfcc",
   474 => x"0c8fde04",
   475 => x"80d1c008",
   476 => x"81e02e09",
   477 => x"81068a38",
   478 => x"810b80cf",
   479 => x"d00c8fde",
   480 => x"0480d1c0",
   481 => x"085280cf",
   482 => x"d008802e",
   483 => x"893880d1",
   484 => x"c0088180",
   485 => x"05527184",
   486 => x"2c728f06",
   487 => x"535380cf",
   488 => x"cc08802e",
   489 => x"9a387284",
   490 => x"2980cf8c",
   491 => x"05721381",
   492 => x"712b7009",
   493 => x"73080673",
   494 => x"0c515353",
   495 => x"8fd20472",
   496 => x"842980cf",
   497 => x"8c057213",
   498 => x"83712b72",
   499 => x"0807720c",
   500 => x"5353800b",
   501 => x"80cfd00c",
   502 => x"800b80cf",
   503 => x"cc0c80d1",
   504 => x"ec5190e5",
   505 => x"2d80d1c0",
   506 => x"08ff24fe",
   507 => x"ea38800b",
   508 => x"80d1c00c",
   509 => x"028c050d",
   510 => x"0402f805",
   511 => x"0d80cf8c",
   512 => x"528f5180",
   513 => x"72708405",
   514 => x"540cff11",
   515 => x"51708025",
   516 => x"f2380288",
   517 => x"050d0402",
   518 => x"f0050d75",
   519 => x"518eca2d",
   520 => x"70822cfc",
   521 => x"0680cf8c",
   522 => x"1172109e",
   523 => x"06710870",
   524 => x"722a7083",
   525 => x"0682742b",
   526 => x"70097406",
   527 => x"760c5451",
   528 => x"56575351",
   529 => x"538ec42d",
   530 => x"7180d1c0",
   531 => x"0c029005",
   532 => x"0d0402fc",
   533 => x"050d7251",
   534 => x"80710c80",
   535 => x"0b84120c",
   536 => x"0284050d",
   537 => x"0402f005",
   538 => x"0d757008",
   539 => x"84120853",
   540 => x"5353ff54",
   541 => x"71712ea8",
   542 => x"388eca2d",
   543 => x"84130870",
   544 => x"84291488",
   545 => x"11700870",
   546 => x"81ff0684",
   547 => x"18088111",
   548 => x"8706841a",
   549 => x"0c535155",
   550 => x"5151518e",
   551 => x"c42d7154",
   552 => x"7380d1c0",
   553 => x"0c029005",
   554 => x"0d0402f4",
   555 => x"050d8eca",
   556 => x"2de00870",
   557 => x"8b2a7081",
   558 => x"06515253",
   559 => x"70802ea1",
   560 => x"3880d1ec",
   561 => x"08708429",
   562 => x"80d1f405",
   563 => x"7481ff06",
   564 => x"710c5151",
   565 => x"80d1ec08",
   566 => x"81118706",
   567 => x"80d1ec0c",
   568 => x"51728c2c",
   569 => x"83ff0680",
   570 => x"d2940c80",
   571 => x"0b80d298",
   572 => x"0c8ebc2d",
   573 => x"8ec42d02",
   574 => x"8c050d04",
   575 => x"02fc050d",
   576 => x"8eca2d81",
   577 => x"0b80d298",
   578 => x"0c8ec42d",
   579 => x"80d29808",
   580 => x"5170f938",
   581 => x"0284050d",
   582 => x"0402fc05",
   583 => x"0d80d1ec",
   584 => x"5190d22d",
   585 => x"8ff92d91",
   586 => x"aa518eb8",
   587 => x"2d028405",
   588 => x"0d0402fc",
   589 => x"050d8fcf",
   590 => x"5186ec2d",
   591 => x"ff115170",
   592 => x"8025f638",
   593 => x"0284050d",
   594 => x"0480d2a0",
   595 => x"0880d1c0",
   596 => x"0c0402fc",
   597 => x"050d810b",
   598 => x"80d0800c",
   599 => x"8151858d",
   600 => x"2d028405",
   601 => x"0d0402fc",
   602 => x"050d92f0",
   603 => x"048ed02d",
   604 => x"80f65190",
   605 => x"972d80d1",
   606 => x"c008f238",
   607 => x"80da5190",
   608 => x"972d80d1",
   609 => x"c008e638",
   610 => x"80cffc08",
   611 => x"5190972d",
   612 => x"80d1c008",
   613 => x"d83880d1",
   614 => x"c00880d0",
   615 => x"800c80d1",
   616 => x"c0085185",
   617 => x"8d2d0284",
   618 => x"050d0402",
   619 => x"ec050d76",
   620 => x"54805287",
   621 => x"0b881580",
   622 => x"f52d5653",
   623 => x"74722483",
   624 => x"38a05372",
   625 => x"5183842d",
   626 => x"81128b15",
   627 => x"80f52d54",
   628 => x"52727225",
   629 => x"de380294",
   630 => x"050d0402",
   631 => x"f0050d80",
   632 => x"d2a00854",
   633 => x"81f92d80",
   634 => x"0b80d2a4",
   635 => x"0c730880",
   636 => x"2e818938",
   637 => x"820b80d1",
   638 => x"d40c80d2",
   639 => x"a4088f06",
   640 => x"80d1d00c",
   641 => x"73085271",
   642 => x"832e9638",
   643 => x"71832689",
   644 => x"3871812e",
   645 => x"b03894e5",
   646 => x"0471852e",
   647 => x"a03894e5",
   648 => x"04881480",
   649 => x"f52d8415",
   650 => x"0880c7c4",
   651 => x"53545286",
   652 => x"c52d7184",
   653 => x"29137008",
   654 => x"525294e9",
   655 => x"04735193",
   656 => x"ab2d94e5",
   657 => x"0480cfd4",
   658 => x"08881508",
   659 => x"2c708106",
   660 => x"51527180",
   661 => x"2e883880",
   662 => x"c7c85194",
   663 => x"e20480c7",
   664 => x"cc5186c5",
   665 => x"2d841408",
   666 => x"5186c52d",
   667 => x"80d2a408",
   668 => x"810580d2",
   669 => x"a40c8c14",
   670 => x"5493ed04",
   671 => x"0290050d",
   672 => x"047180d2",
   673 => x"a00c93db",
   674 => x"2d80d2a4",
   675 => x"08ff0580",
   676 => x"d2a80c04",
   677 => x"02e8050d",
   678 => x"80d2a008",
   679 => x"80d2ac08",
   680 => x"575580f6",
   681 => x"5190972d",
   682 => x"80d1c008",
   683 => x"812a7081",
   684 => x"06515271",
   685 => x"802ea238",
   686 => x"95be048e",
   687 => x"d02d80f6",
   688 => x"5190972d",
   689 => x"80d1c008",
   690 => x"f23880d0",
   691 => x"80088132",
   692 => x"7080d080",
   693 => x"0c51858d",
   694 => x"2d800b80",
   695 => x"d29c0c86",
   696 => x"5190972d",
   697 => x"80d1c008",
   698 => x"812a7081",
   699 => x"06515271",
   700 => x"802e8b38",
   701 => x"80c98008",
   702 => x"903280c9",
   703 => x"800c8c51",
   704 => x"90972d80",
   705 => x"d1c00881",
   706 => x"2a708106",
   707 => x"51527180",
   708 => x"2e80d138",
   709 => x"80cfd808",
   710 => x"80cfec08",
   711 => x"80cfd80c",
   712 => x"80cfec0c",
   713 => x"80cfdc08",
   714 => x"80cff008",
   715 => x"80cfdc0c",
   716 => x"80cff00c",
   717 => x"80cfe008",
   718 => x"80cff408",
   719 => x"80cfe00c",
   720 => x"80cff40c",
   721 => x"80cfe408",
   722 => x"80cff808",
   723 => x"80cfe40c",
   724 => x"80cff80c",
   725 => x"80cfe808",
   726 => x"80cffc08",
   727 => x"80cfe80c",
   728 => x"80cffc0c",
   729 => x"80d29408",
   730 => x"a0065280",
   731 => x"72259638",
   732 => x"92b22d8e",
   733 => x"d02d80d0",
   734 => x"80088132",
   735 => x"7080d080",
   736 => x"0c51858d",
   737 => x"2d80d080",
   738 => x"0882ef38",
   739 => x"80cfec08",
   740 => x"5190972d",
   741 => x"80d1c008",
   742 => x"802e8b38",
   743 => x"80d29c08",
   744 => x"810780d2",
   745 => x"9c0c80cf",
   746 => x"f0085190",
   747 => x"972d80d1",
   748 => x"c008802e",
   749 => x"8b3880d2",
   750 => x"9c088207",
   751 => x"80d29c0c",
   752 => x"80cff408",
   753 => x"5190972d",
   754 => x"80d1c008",
   755 => x"802e8b38",
   756 => x"80d29c08",
   757 => x"840780d2",
   758 => x"9c0c80cf",
   759 => x"f8085190",
   760 => x"972d80d1",
   761 => x"c008802e",
   762 => x"8b3880d2",
   763 => x"9c088807",
   764 => x"80d29c0c",
   765 => x"80cffc08",
   766 => x"5190972d",
   767 => x"80d1c008",
   768 => x"802e8b38",
   769 => x"80d29c08",
   770 => x"900780d2",
   771 => x"9c0c80cf",
   772 => x"d8085190",
   773 => x"972d80d1",
   774 => x"c008802e",
   775 => x"8c3880d2",
   776 => x"9c088280",
   777 => x"0780d29c",
   778 => x"0c80cfdc",
   779 => x"08519097",
   780 => x"2d80d1c0",
   781 => x"08802e8c",
   782 => x"3880d29c",
   783 => x"08848007",
   784 => x"80d29c0c",
   785 => x"80cfe008",
   786 => x"5190972d",
   787 => x"80d1c008",
   788 => x"802e8c38",
   789 => x"80d29c08",
   790 => x"88800780",
   791 => x"d29c0c80",
   792 => x"cfe40851",
   793 => x"90972d80",
   794 => x"d1c00880",
   795 => x"2e8c3880",
   796 => x"d29c0890",
   797 => x"800780d2",
   798 => x"9c0c80cf",
   799 => x"e8085190",
   800 => x"972d80d1",
   801 => x"c008802e",
   802 => x"8c3880d2",
   803 => x"9c08a080",
   804 => x"0780d29c",
   805 => x"0c945190",
   806 => x"972d80d1",
   807 => x"c0085291",
   808 => x"5190972d",
   809 => x"7180d1c0",
   810 => x"08065280",
   811 => x"e6519097",
   812 => x"2d7180d1",
   813 => x"c0080652",
   814 => x"71802e8d",
   815 => x"3880d29c",
   816 => x"08848080",
   817 => x"0780d29c",
   818 => x"0c80fe51",
   819 => x"90972d80",
   820 => x"d1c00852",
   821 => x"87519097",
   822 => x"2d7180d1",
   823 => x"c0080752",
   824 => x"71802e8d",
   825 => x"3880d29c",
   826 => x"08888080",
   827 => x"0780d29c",
   828 => x"0c80d29c",
   829 => x"08ed0ca2",
   830 => x"85049451",
   831 => x"90972d80",
   832 => x"d1c00852",
   833 => x"91519097",
   834 => x"2d7180d1",
   835 => x"c0080652",
   836 => x"80e65190",
   837 => x"972d7180",
   838 => x"d1c00806",
   839 => x"5271802e",
   840 => x"8d3880d2",
   841 => x"9c088480",
   842 => x"800780d2",
   843 => x"9c0c80fe",
   844 => x"5190972d",
   845 => x"80d1c008",
   846 => x"52875190",
   847 => x"972d7180",
   848 => x"d1c00807",
   849 => x"5271802e",
   850 => x"8d3880d2",
   851 => x"9c088880",
   852 => x"800780d2",
   853 => x"9c0c80d2",
   854 => x"9c08ed0c",
   855 => x"81f55190",
   856 => x"972d80d1",
   857 => x"c008812a",
   858 => x"70810651",
   859 => x"5271a438",
   860 => x"80cfec08",
   861 => x"5190972d",
   862 => x"80d1c008",
   863 => x"812a7081",
   864 => x"06515271",
   865 => x"8e3880d2",
   866 => x"94088106",
   867 => x"52807225",
   868 => x"80c23880",
   869 => x"d2940881",
   870 => x"06528072",
   871 => x"25843892",
   872 => x"b22d80d2",
   873 => x"a8085271",
   874 => x"802e8a38",
   875 => x"ff1280d2",
   876 => x"a80c9bd4",
   877 => x"0480d2a4",
   878 => x"081080d2",
   879 => x"a4080570",
   880 => x"84291651",
   881 => x"52881208",
   882 => x"802e8938",
   883 => x"ff518812",
   884 => x"0852712d",
   885 => x"81f25190",
   886 => x"972d80d1",
   887 => x"c008812a",
   888 => x"70810651",
   889 => x"5271a438",
   890 => x"80cff008",
   891 => x"5190972d",
   892 => x"80d1c008",
   893 => x"812a7081",
   894 => x"06515271",
   895 => x"8e3880d2",
   896 => x"94088206",
   897 => x"52807225",
   898 => x"80c33880",
   899 => x"d2940882",
   900 => x"06528072",
   901 => x"25843892",
   902 => x"b22d80d2",
   903 => x"a408ff11",
   904 => x"80d2a808",
   905 => x"56535373",
   906 => x"72258a38",
   907 => x"811480d2",
   908 => x"a80c9ccd",
   909 => x"04721013",
   910 => x"70842916",
   911 => x"51528812",
   912 => x"08802e89",
   913 => x"38fe5188",
   914 => x"12085271",
   915 => x"2d81fd51",
   916 => x"90972d80",
   917 => x"d1c00881",
   918 => x"2a708106",
   919 => x"515271a4",
   920 => x"3880cff4",
   921 => x"08519097",
   922 => x"2d80d1c0",
   923 => x"08812a70",
   924 => x"81065152",
   925 => x"718e3880",
   926 => x"d2940884",
   927 => x"06528072",
   928 => x"2580c038",
   929 => x"80d29408",
   930 => x"84065280",
   931 => x"72258438",
   932 => x"92b22d80",
   933 => x"d2a80880",
   934 => x"2e8a3880",
   935 => x"0b80d2a8",
   936 => x"0c9dc304",
   937 => x"80d2a408",
   938 => x"1080d2a4",
   939 => x"08057084",
   940 => x"29165152",
   941 => x"88120880",
   942 => x"2e8938fd",
   943 => x"51881208",
   944 => x"52712d81",
   945 => x"fa519097",
   946 => x"2d80d1c0",
   947 => x"08812a70",
   948 => x"81065152",
   949 => x"71a43880",
   950 => x"cff80851",
   951 => x"90972d80",
   952 => x"d1c00881",
   953 => x"2a708106",
   954 => x"5152718e",
   955 => x"3880d294",
   956 => x"08880652",
   957 => x"80722580",
   958 => x"c03880d2",
   959 => x"94088806",
   960 => x"52807225",
   961 => x"843892b2",
   962 => x"2d80d2a4",
   963 => x"08ff1154",
   964 => x"5280d2a8",
   965 => x"08732589",
   966 => x"387280d2",
   967 => x"a80c9eb9",
   968 => x"04711012",
   969 => x"70842916",
   970 => x"51528812",
   971 => x"08802e89",
   972 => x"38fc5188",
   973 => x"12085271",
   974 => x"2d80d2a8",
   975 => x"08705354",
   976 => x"73802e8a",
   977 => x"388c15ff",
   978 => x"1555559e",
   979 => x"c004820b",
   980 => x"80d1d40c",
   981 => x"718f0680",
   982 => x"d1d00c81",
   983 => x"eb519097",
   984 => x"2d80d1c0",
   985 => x"08812a70",
   986 => x"81065152",
   987 => x"71802ead",
   988 => x"38740885",
   989 => x"2e098106",
   990 => x"a4388815",
   991 => x"80f52dff",
   992 => x"05527188",
   993 => x"1681b72d",
   994 => x"71982b52",
   995 => x"71802588",
   996 => x"38800b88",
   997 => x"1681b72d",
   998 => x"745193ab",
   999 => x"2d81f451",
  1000 => x"90972d80",
  1001 => x"d1c00881",
  1002 => x"2a708106",
  1003 => x"51527180",
  1004 => x"2eb33874",
  1005 => x"08852e09",
  1006 => x"8106aa38",
  1007 => x"881580f5",
  1008 => x"2d810552",
  1009 => x"71881681",
  1010 => x"b72d7181",
  1011 => x"ff068b16",
  1012 => x"80f52d54",
  1013 => x"52727227",
  1014 => x"87387288",
  1015 => x"1681b72d",
  1016 => x"745193ab",
  1017 => x"2d80da51",
  1018 => x"90972d80",
  1019 => x"d1c00881",
  1020 => x"2a708106",
  1021 => x"5152718e",
  1022 => x"3880d294",
  1023 => x"08900652",
  1024 => x"80722581",
  1025 => x"bc3880d2",
  1026 => x"a00880d2",
  1027 => x"94089006",
  1028 => x"53538072",
  1029 => x"25843892",
  1030 => x"b22d80d2",
  1031 => x"a8085473",
  1032 => x"802e8a38",
  1033 => x"8c13ff15",
  1034 => x"5553a09f",
  1035 => x"04720852",
  1036 => x"71822ea6",
  1037 => x"38718226",
  1038 => x"89387181",
  1039 => x"2eaa38a1",
  1040 => x"c1047183",
  1041 => x"2eb43871",
  1042 => x"842e0981",
  1043 => x"0680f238",
  1044 => x"88130851",
  1045 => x"95812da1",
  1046 => x"c10480d2",
  1047 => x"a8085188",
  1048 => x"13085271",
  1049 => x"2da1c104",
  1050 => x"810b8814",
  1051 => x"082b80cf",
  1052 => x"d4083280",
  1053 => x"cfd40ca1",
  1054 => x"95048813",
  1055 => x"80f52d81",
  1056 => x"058b1480",
  1057 => x"f52d5354",
  1058 => x"71742483",
  1059 => x"38805473",
  1060 => x"881481b7",
  1061 => x"2d93db2d",
  1062 => x"a1c10475",
  1063 => x"08802ea4",
  1064 => x"38750851",
  1065 => x"90972d80",
  1066 => x"d1c00881",
  1067 => x"06527180",
  1068 => x"2e8c3880",
  1069 => x"d2a80851",
  1070 => x"84160852",
  1071 => x"712d8816",
  1072 => x"5675d838",
  1073 => x"8054800b",
  1074 => x"80d1d40c",
  1075 => x"738f0680",
  1076 => x"d1d00ca0",
  1077 => x"527380d2",
  1078 => x"a8082e09",
  1079 => x"81069938",
  1080 => x"80d2a408",
  1081 => x"ff057432",
  1082 => x"70098105",
  1083 => x"7072079f",
  1084 => x"2a917131",
  1085 => x"51515353",
  1086 => x"71518384",
  1087 => x"2d811454",
  1088 => x"8e7425c2",
  1089 => x"3880d080",
  1090 => x"0880d1c0",
  1091 => x"0c029805",
  1092 => x"0d0402f4",
  1093 => x"050dd452",
  1094 => x"81ff720c",
  1095 => x"71085381",
  1096 => x"ff720c72",
  1097 => x"882b83fe",
  1098 => x"80067208",
  1099 => x"7081ff06",
  1100 => x"51525381",
  1101 => x"ff720c72",
  1102 => x"7107882b",
  1103 => x"72087081",
  1104 => x"ff065152",
  1105 => x"5381ff72",
  1106 => x"0c727107",
  1107 => x"882b7208",
  1108 => x"7081ff06",
  1109 => x"720780d1",
  1110 => x"c00c5253",
  1111 => x"028c050d",
  1112 => x"0402f405",
  1113 => x"0d747671",
  1114 => x"81ff06d4",
  1115 => x"0c535380",
  1116 => x"d2b00885",
  1117 => x"3871892b",
  1118 => x"5271982a",
  1119 => x"d40c7190",
  1120 => x"2a7081ff",
  1121 => x"06d40c51",
  1122 => x"71882a70",
  1123 => x"81ff06d4",
  1124 => x"0c517181",
  1125 => x"ff06d40c",
  1126 => x"72902a70",
  1127 => x"81ff06d4",
  1128 => x"0c51d408",
  1129 => x"7081ff06",
  1130 => x"515182b8",
  1131 => x"bf527081",
  1132 => x"ff2e0981",
  1133 => x"06943881",
  1134 => x"ff0bd40c",
  1135 => x"d4087081",
  1136 => x"ff06ff14",
  1137 => x"54515171",
  1138 => x"e5387080",
  1139 => x"d1c00c02",
  1140 => x"8c050d04",
  1141 => x"02fc050d",
  1142 => x"81c75181",
  1143 => x"ff0bd40c",
  1144 => x"ff115170",
  1145 => x"8025f438",
  1146 => x"0284050d",
  1147 => x"0402f405",
  1148 => x"0d81ff0b",
  1149 => x"d40c9353",
  1150 => x"805287fc",
  1151 => x"80c151a2",
  1152 => x"e12d80d1",
  1153 => x"c0088b38",
  1154 => x"81ff0bd4",
  1155 => x"0c8153a4",
  1156 => x"9b04a3d4",
  1157 => x"2dff1353",
  1158 => x"72de3872",
  1159 => x"80d1c00c",
  1160 => x"028c050d",
  1161 => x"0402ec05",
  1162 => x"0d810b80",
  1163 => x"d2b00c84",
  1164 => x"54d00870",
  1165 => x"8f2a7081",
  1166 => x"06515153",
  1167 => x"72f33872",
  1168 => x"d00ca3d4",
  1169 => x"2d80c7d0",
  1170 => x"5186c52d",
  1171 => x"d008708f",
  1172 => x"2a708106",
  1173 => x"51515372",
  1174 => x"f338810b",
  1175 => x"d00cb153",
  1176 => x"805284d4",
  1177 => x"80c051a2",
  1178 => x"e12d80d1",
  1179 => x"c008812e",
  1180 => x"93387282",
  1181 => x"2ebf38ff",
  1182 => x"135372e4",
  1183 => x"38ff1454",
  1184 => x"73ffae38",
  1185 => x"a3d42d83",
  1186 => x"aa52849c",
  1187 => x"80c851a2",
  1188 => x"e12d80d1",
  1189 => x"c008812e",
  1190 => x"09810693",
  1191 => x"38a2922d",
  1192 => x"80d1c008",
  1193 => x"83ffff06",
  1194 => x"537283aa",
  1195 => x"2e9f38a3",
  1196 => x"ed2da5c8",
  1197 => x"0480c7dc",
  1198 => x"5186c52d",
  1199 => x"8053a79d",
  1200 => x"0480c7f4",
  1201 => x"5186c52d",
  1202 => x"8054a6ee",
  1203 => x"0481ff0b",
  1204 => x"d40cb154",
  1205 => x"a3d42d8f",
  1206 => x"cf538052",
  1207 => x"87fc80f7",
  1208 => x"51a2e12d",
  1209 => x"80d1c008",
  1210 => x"5580d1c0",
  1211 => x"08812e09",
  1212 => x"81069c38",
  1213 => x"81ff0bd4",
  1214 => x"0c820a52",
  1215 => x"849c80e9",
  1216 => x"51a2e12d",
  1217 => x"80d1c008",
  1218 => x"802e8d38",
  1219 => x"a3d42dff",
  1220 => x"135372c6",
  1221 => x"38a6e104",
  1222 => x"81ff0bd4",
  1223 => x"0c80d1c0",
  1224 => x"085287fc",
  1225 => x"80fa51a2",
  1226 => x"e12d80d1",
  1227 => x"c008b238",
  1228 => x"81ff0bd4",
  1229 => x"0cd40853",
  1230 => x"81ff0bd4",
  1231 => x"0c81ff0b",
  1232 => x"d40c81ff",
  1233 => x"0bd40c81",
  1234 => x"ff0bd40c",
  1235 => x"72862a70",
  1236 => x"81067656",
  1237 => x"51537296",
  1238 => x"3880d1c0",
  1239 => x"0854a6ee",
  1240 => x"0473822e",
  1241 => x"fedb38ff",
  1242 => x"145473fe",
  1243 => x"e7387380",
  1244 => x"d2b00c73",
  1245 => x"8b388152",
  1246 => x"87fc80d0",
  1247 => x"51a2e12d",
  1248 => x"81ff0bd4",
  1249 => x"0cd00870",
  1250 => x"8f2a7081",
  1251 => x"06515153",
  1252 => x"72f33872",
  1253 => x"d00c81ff",
  1254 => x"0bd40c81",
  1255 => x"537280d1",
  1256 => x"c00c0294",
  1257 => x"050d0402",
  1258 => x"e8050d78",
  1259 => x"55805681",
  1260 => x"ff0bd40c",
  1261 => x"d008708f",
  1262 => x"2a708106",
  1263 => x"51515372",
  1264 => x"f3388281",
  1265 => x"0bd00c81",
  1266 => x"ff0bd40c",
  1267 => x"775287fc",
  1268 => x"80d151a2",
  1269 => x"e12d80db",
  1270 => x"c6df5480",
  1271 => x"d1c00880",
  1272 => x"2e8b3880",
  1273 => x"c8945186",
  1274 => x"c52da8c1",
  1275 => x"0481ff0b",
  1276 => x"d40cd408",
  1277 => x"7081ff06",
  1278 => x"51537281",
  1279 => x"fe2e0981",
  1280 => x"069e3880",
  1281 => x"ff53a292",
  1282 => x"2d80d1c0",
  1283 => x"08757084",
  1284 => x"05570cff",
  1285 => x"13537280",
  1286 => x"25ec3881",
  1287 => x"56a8a604",
  1288 => x"ff145473",
  1289 => x"c83881ff",
  1290 => x"0bd40c81",
  1291 => x"ff0bd40c",
  1292 => x"d008708f",
  1293 => x"2a708106",
  1294 => x"51515372",
  1295 => x"f33872d0",
  1296 => x"0c7580d1",
  1297 => x"c00c0298",
  1298 => x"050d0402",
  1299 => x"e8050d77",
  1300 => x"797b5855",
  1301 => x"55805372",
  1302 => x"7625a338",
  1303 => x"74708105",
  1304 => x"5680f52d",
  1305 => x"74708105",
  1306 => x"5680f52d",
  1307 => x"52527171",
  1308 => x"2e863881",
  1309 => x"51a98004",
  1310 => x"811353a8",
  1311 => x"d7048051",
  1312 => x"7080d1c0",
  1313 => x"0c029805",
  1314 => x"0d0402ec",
  1315 => x"050d7655",
  1316 => x"74802e80",
  1317 => x"c2389a15",
  1318 => x"80e02d51",
  1319 => x"b79f2d80",
  1320 => x"d1c00880",
  1321 => x"d1c00880",
  1322 => x"d8e40c80",
  1323 => x"d1c00854",
  1324 => x"5480d8c0",
  1325 => x"08802e9a",
  1326 => x"38941580",
  1327 => x"e02d51b7",
  1328 => x"9f2d80d1",
  1329 => x"c008902b",
  1330 => x"83fff00a",
  1331 => x"06707507",
  1332 => x"51537280",
  1333 => x"d8e40c80",
  1334 => x"d8e40853",
  1335 => x"72802e9d",
  1336 => x"3880d8b8",
  1337 => x"08fe1471",
  1338 => x"2980d8cc",
  1339 => x"080580d8",
  1340 => x"e80c7084",
  1341 => x"2b80d8c4",
  1342 => x"0c54aaab",
  1343 => x"0480d8d0",
  1344 => x"0880d8e4",
  1345 => x"0c80d8d4",
  1346 => x"0880d8e8",
  1347 => x"0c80d8c0",
  1348 => x"08802e8b",
  1349 => x"3880d8b8",
  1350 => x"08842b53",
  1351 => x"aaa60480",
  1352 => x"d8d80884",
  1353 => x"2b537280",
  1354 => x"d8c40c02",
  1355 => x"94050d04",
  1356 => x"02d8050d",
  1357 => x"800b80d8",
  1358 => x"c00c8454",
  1359 => x"a4a52d80",
  1360 => x"d1c00880",
  1361 => x"2e973880",
  1362 => x"d2b45280",
  1363 => x"51a7a72d",
  1364 => x"80d1c008",
  1365 => x"802e8638",
  1366 => x"fe54aae5",
  1367 => x"04ff1454",
  1368 => x"738024d8",
  1369 => x"38738d38",
  1370 => x"80c8a451",
  1371 => x"86c52d73",
  1372 => x"55b0ba04",
  1373 => x"8056810b",
  1374 => x"80d8ec0c",
  1375 => x"885380c8",
  1376 => x"b85280d2",
  1377 => x"ea51a8cb",
  1378 => x"2d80d1c0",
  1379 => x"08762e09",
  1380 => x"81068938",
  1381 => x"80d1c008",
  1382 => x"80d8ec0c",
  1383 => x"885380c8",
  1384 => x"c45280d3",
  1385 => x"8651a8cb",
  1386 => x"2d80d1c0",
  1387 => x"08893880",
  1388 => x"d1c00880",
  1389 => x"d8ec0c80",
  1390 => x"d8ec0880",
  1391 => x"2e818138",
  1392 => x"80d5fa0b",
  1393 => x"80f52d80",
  1394 => x"d5fb0b80",
  1395 => x"f52d7198",
  1396 => x"2b71902b",
  1397 => x"0780d5fc",
  1398 => x"0b80f52d",
  1399 => x"70882b72",
  1400 => x"0780d5fd",
  1401 => x"0b80f52d",
  1402 => x"710780d6",
  1403 => x"b20b80f5",
  1404 => x"2d80d6b3",
  1405 => x"0b80f52d",
  1406 => x"71882b07",
  1407 => x"535f5452",
  1408 => x"5a565755",
  1409 => x"7381abaa",
  1410 => x"2e098106",
  1411 => x"8e387551",
  1412 => x"b6ee2d80",
  1413 => x"d1c00856",
  1414 => x"aca90473",
  1415 => x"82d4d52e",
  1416 => x"883880c8",
  1417 => x"d051acf5",
  1418 => x"0480d2b4",
  1419 => x"527551a7",
  1420 => x"a72d80d1",
  1421 => x"c0085580",
  1422 => x"d1c00880",
  1423 => x"2e83fb38",
  1424 => x"885380c8",
  1425 => x"c45280d3",
  1426 => x"8651a8cb",
  1427 => x"2d80d1c0",
  1428 => x"088a3881",
  1429 => x"0b80d8c0",
  1430 => x"0cacfb04",
  1431 => x"885380c8",
  1432 => x"b85280d2",
  1433 => x"ea51a8cb",
  1434 => x"2d80d1c0",
  1435 => x"08802e8b",
  1436 => x"3880c8e4",
  1437 => x"5186c52d",
  1438 => x"adda0480",
  1439 => x"d6b20b80",
  1440 => x"f52d5473",
  1441 => x"80d52e09",
  1442 => x"810680ce",
  1443 => x"3880d6b3",
  1444 => x"0b80f52d",
  1445 => x"547381aa",
  1446 => x"2e098106",
  1447 => x"bd38800b",
  1448 => x"80d2b40b",
  1449 => x"80f52d56",
  1450 => x"547481e9",
  1451 => x"2e833881",
  1452 => x"547481eb",
  1453 => x"2e8c3880",
  1454 => x"5573752e",
  1455 => x"09810682",
  1456 => x"f93880d2",
  1457 => x"bf0b80f5",
  1458 => x"2d55748e",
  1459 => x"3880d2c0",
  1460 => x"0b80f52d",
  1461 => x"5473822e",
  1462 => x"86388055",
  1463 => x"b0ba0480",
  1464 => x"d2c10b80",
  1465 => x"f52d7080",
  1466 => x"d8b80cff",
  1467 => x"0580d8bc",
  1468 => x"0c80d2c2",
  1469 => x"0b80f52d",
  1470 => x"80d2c30b",
  1471 => x"80f52d58",
  1472 => x"76057782",
  1473 => x"80290570",
  1474 => x"80d8c80c",
  1475 => x"80d2c40b",
  1476 => x"80f52d70",
  1477 => x"80d8dc0c",
  1478 => x"80d8c008",
  1479 => x"59575876",
  1480 => x"802e81b7",
  1481 => x"38885380",
  1482 => x"c8c45280",
  1483 => x"d38651a8",
  1484 => x"cb2d80d1",
  1485 => x"c0088282",
  1486 => x"3880d8b8",
  1487 => x"0870842b",
  1488 => x"80d8c40c",
  1489 => x"7080d8d8",
  1490 => x"0c80d2d9",
  1491 => x"0b80f52d",
  1492 => x"80d2d80b",
  1493 => x"80f52d71",
  1494 => x"82802905",
  1495 => x"80d2da0b",
  1496 => x"80f52d70",
  1497 => x"84808029",
  1498 => x"1280d2db",
  1499 => x"0b80f52d",
  1500 => x"7081800a",
  1501 => x"29127080",
  1502 => x"d8e00c80",
  1503 => x"d8dc0871",
  1504 => x"2980d8c8",
  1505 => x"08057080",
  1506 => x"d8cc0c80",
  1507 => x"d2e10b80",
  1508 => x"f52d80d2",
  1509 => x"e00b80f5",
  1510 => x"2d718280",
  1511 => x"290580d2",
  1512 => x"e20b80f5",
  1513 => x"2d708480",
  1514 => x"80291280",
  1515 => x"d2e30b80",
  1516 => x"f52d7098",
  1517 => x"2b81f00a",
  1518 => x"06720570",
  1519 => x"80d8d00c",
  1520 => x"fe117e29",
  1521 => x"770580d8",
  1522 => x"d40c5259",
  1523 => x"5243545e",
  1524 => x"51525952",
  1525 => x"5d575957",
  1526 => x"b0b30480",
  1527 => x"d2c60b80",
  1528 => x"f52d80d2",
  1529 => x"c50b80f5",
  1530 => x"2d718280",
  1531 => x"29057080",
  1532 => x"d8c40c70",
  1533 => x"a02983ff",
  1534 => x"0570892a",
  1535 => x"7080d8d8",
  1536 => x"0c80d2cb",
  1537 => x"0b80f52d",
  1538 => x"80d2ca0b",
  1539 => x"80f52d71",
  1540 => x"82802905",
  1541 => x"7080d8e0",
  1542 => x"0c7b7129",
  1543 => x"1e7080d8",
  1544 => x"d40c7d80",
  1545 => x"d8d00c73",
  1546 => x"0580d8cc",
  1547 => x"0c555e51",
  1548 => x"51555580",
  1549 => x"51a98a2d",
  1550 => x"81557480",
  1551 => x"d1c00c02",
  1552 => x"a8050d04",
  1553 => x"02ec050d",
  1554 => x"7670872c",
  1555 => x"7180ff06",
  1556 => x"55565480",
  1557 => x"d8c0088a",
  1558 => x"3873882c",
  1559 => x"7481ff06",
  1560 => x"545580d2",
  1561 => x"b45280d8",
  1562 => x"c8081551",
  1563 => x"a7a72d80",
  1564 => x"d1c00854",
  1565 => x"80d1c008",
  1566 => x"802eb838",
  1567 => x"80d8c008",
  1568 => x"802e9a38",
  1569 => x"72842980",
  1570 => x"d2b40570",
  1571 => x"085253b6",
  1572 => x"ee2d80d1",
  1573 => x"c008f00a",
  1574 => x"0653b1b1",
  1575 => x"04721080",
  1576 => x"d2b40570",
  1577 => x"80e02d52",
  1578 => x"53b79f2d",
  1579 => x"80d1c008",
  1580 => x"53725473",
  1581 => x"80d1c00c",
  1582 => x"0294050d",
  1583 => x"0402e005",
  1584 => x"0d797084",
  1585 => x"2c80d8e8",
  1586 => x"0805718f",
  1587 => x"06525553",
  1588 => x"728a3880",
  1589 => x"d2b45273",
  1590 => x"51a7a72d",
  1591 => x"72a02980",
  1592 => x"d2b40554",
  1593 => x"807480f5",
  1594 => x"2d565374",
  1595 => x"732e8338",
  1596 => x"81537481",
  1597 => x"e52e81f4",
  1598 => x"38817074",
  1599 => x"06545872",
  1600 => x"802e81e8",
  1601 => x"388b1480",
  1602 => x"f52d7083",
  1603 => x"2a790658",
  1604 => x"56769b38",
  1605 => x"80d08408",
  1606 => x"53728938",
  1607 => x"7280d6b4",
  1608 => x"0b81b72d",
  1609 => x"7680d084",
  1610 => x"0c7353b3",
  1611 => x"ee04758f",
  1612 => x"2e098106",
  1613 => x"81b63874",
  1614 => x"9f068d29",
  1615 => x"80d6a711",
  1616 => x"51538114",
  1617 => x"80f52d73",
  1618 => x"70810555",
  1619 => x"81b72d83",
  1620 => x"1480f52d",
  1621 => x"73708105",
  1622 => x"5581b72d",
  1623 => x"851480f5",
  1624 => x"2d737081",
  1625 => x"055581b7",
  1626 => x"2d871480",
  1627 => x"f52d7370",
  1628 => x"81055581",
  1629 => x"b72d8914",
  1630 => x"80f52d73",
  1631 => x"70810555",
  1632 => x"81b72d8e",
  1633 => x"1480f52d",
  1634 => x"73708105",
  1635 => x"5581b72d",
  1636 => x"901480f5",
  1637 => x"2d737081",
  1638 => x"055581b7",
  1639 => x"2d921480",
  1640 => x"f52d7370",
  1641 => x"81055581",
  1642 => x"b72d9414",
  1643 => x"80f52d73",
  1644 => x"70810555",
  1645 => x"81b72d96",
  1646 => x"1480f52d",
  1647 => x"73708105",
  1648 => x"5581b72d",
  1649 => x"981480f5",
  1650 => x"2d737081",
  1651 => x"055581b7",
  1652 => x"2d9c1480",
  1653 => x"f52d7370",
  1654 => x"81055581",
  1655 => x"b72d9e14",
  1656 => x"80f52d73",
  1657 => x"81b72d77",
  1658 => x"80d0840c",
  1659 => x"80537280",
  1660 => x"d1c00c02",
  1661 => x"a0050d04",
  1662 => x"02cc050d",
  1663 => x"7e605e5a",
  1664 => x"800b80d8",
  1665 => x"e40880d8",
  1666 => x"e808595c",
  1667 => x"56805880",
  1668 => x"d8c40878",
  1669 => x"2e81b838",
  1670 => x"778f06a0",
  1671 => x"17575473",
  1672 => x"913880d2",
  1673 => x"b4527651",
  1674 => x"811757a7",
  1675 => x"a72d80d2",
  1676 => x"b4568076",
  1677 => x"80f52d56",
  1678 => x"5474742e",
  1679 => x"83388154",
  1680 => x"7481e52e",
  1681 => x"80fd3881",
  1682 => x"70750655",
  1683 => x"5c73802e",
  1684 => x"80f1388b",
  1685 => x"1680f52d",
  1686 => x"98065978",
  1687 => x"80e5388b",
  1688 => x"537c5275",
  1689 => x"51a8cb2d",
  1690 => x"80d1c008",
  1691 => x"80d5389c",
  1692 => x"160851b6",
  1693 => x"ee2d80d1",
  1694 => x"c008841b",
  1695 => x"0c9a1680",
  1696 => x"e02d51b7",
  1697 => x"9f2d80d1",
  1698 => x"c00880d1",
  1699 => x"c008881c",
  1700 => x"0c80d1c0",
  1701 => x"08555580",
  1702 => x"d8c00880",
  1703 => x"2e993894",
  1704 => x"1680e02d",
  1705 => x"51b79f2d",
  1706 => x"80d1c008",
  1707 => x"902b83ff",
  1708 => x"f00a0670",
  1709 => x"16515473",
  1710 => x"881b0c78",
  1711 => x"7a0c7b54",
  1712 => x"b68b0481",
  1713 => x"185880d8",
  1714 => x"c4087826",
  1715 => x"feca3880",
  1716 => x"d8c00880",
  1717 => x"2eb3387a",
  1718 => x"51b0c42d",
  1719 => x"80d1c008",
  1720 => x"80d1c008",
  1721 => x"80ffffff",
  1722 => x"f806555b",
  1723 => x"7380ffff",
  1724 => x"fff82e95",
  1725 => x"3880d1c0",
  1726 => x"08fe0580",
  1727 => x"d8b80829",
  1728 => x"80d8cc08",
  1729 => x"0557b48d",
  1730 => x"04805473",
  1731 => x"80d1c00c",
  1732 => x"02b4050d",
  1733 => x"0402f405",
  1734 => x"0d747008",
  1735 => x"8105710c",
  1736 => x"700880d8",
  1737 => x"bc080653",
  1738 => x"53718f38",
  1739 => x"88130851",
  1740 => x"b0c42d80",
  1741 => x"d1c00888",
  1742 => x"140c810b",
  1743 => x"80d1c00c",
  1744 => x"028c050d",
  1745 => x"0402f005",
  1746 => x"0d758811",
  1747 => x"08fe0580",
  1748 => x"d8b80829",
  1749 => x"80d8cc08",
  1750 => x"11720880",
  1751 => x"d8bc0806",
  1752 => x"05795553",
  1753 => x"5454a7a7",
  1754 => x"2d029005",
  1755 => x"0d0402f4",
  1756 => x"050d7470",
  1757 => x"882a83fe",
  1758 => x"80067072",
  1759 => x"982a0772",
  1760 => x"882b87fc",
  1761 => x"80800673",
  1762 => x"982b81f0",
  1763 => x"0a067173",
  1764 => x"070780d1",
  1765 => x"c00c5651",
  1766 => x"5351028c",
  1767 => x"050d0402",
  1768 => x"f8050d02",
  1769 => x"8e0580f5",
  1770 => x"2d74882b",
  1771 => x"077083ff",
  1772 => x"ff0680d1",
  1773 => x"c00c5102",
  1774 => x"88050d04",
  1775 => x"02f4050d",
  1776 => x"74767853",
  1777 => x"54528071",
  1778 => x"25973872",
  1779 => x"70810554",
  1780 => x"80f52d72",
  1781 => x"70810554",
  1782 => x"81b72dff",
  1783 => x"115170eb",
  1784 => x"38807281",
  1785 => x"b72d028c",
  1786 => x"050d0402",
  1787 => x"e8050d77",
  1788 => x"56807056",
  1789 => x"54737624",
  1790 => x"b63880d8",
  1791 => x"c408742e",
  1792 => x"ae387351",
  1793 => x"b1bd2d80",
  1794 => x"d1c00880",
  1795 => x"d1c00809",
  1796 => x"81057080",
  1797 => x"d1c00807",
  1798 => x"9f2a7705",
  1799 => x"81175757",
  1800 => x"53537476",
  1801 => x"24893880",
  1802 => x"d8c40874",
  1803 => x"26d43872",
  1804 => x"80d1c00c",
  1805 => x"0298050d",
  1806 => x"0402ec05",
  1807 => x"0d80d1bc",
  1808 => x"081751b7",
  1809 => x"eb2d80d1",
  1810 => x"c0085580",
  1811 => x"d1c00880",
  1812 => x"2ea2388b",
  1813 => x"5380d1c0",
  1814 => x"085280d6",
  1815 => x"b451b7bc",
  1816 => x"2d80d8f0",
  1817 => x"08547380",
  1818 => x"2e8a3888",
  1819 => x"155280d6",
  1820 => x"b451732d",
  1821 => x"0294050d",
  1822 => x"0402dc05",
  1823 => x"0d80705a",
  1824 => x"557480d1",
  1825 => x"bc0825b4",
  1826 => x"3880d8c4",
  1827 => x"08752eac",
  1828 => x"387851b1",
  1829 => x"bd2d80d1",
  1830 => x"c0080981",
  1831 => x"057080d1",
  1832 => x"c008079f",
  1833 => x"2a760581",
  1834 => x"1b5b5654",
  1835 => x"7480d1bc",
  1836 => x"08258938",
  1837 => x"80d8c408",
  1838 => x"7926d638",
  1839 => x"80557880",
  1840 => x"d8c40827",
  1841 => x"81db3878",
  1842 => x"51b1bd2d",
  1843 => x"80d1c008",
  1844 => x"802e81ad",
  1845 => x"3880d1c0",
  1846 => x"088b0580",
  1847 => x"f52d7084",
  1848 => x"2a708106",
  1849 => x"77107884",
  1850 => x"2b80d6b4",
  1851 => x"0b80f52d",
  1852 => x"5c5c5351",
  1853 => x"55567380",
  1854 => x"2e80cb38",
  1855 => x"7416822b",
  1856 => x"bbc50b80",
  1857 => x"d090120c",
  1858 => x"54777531",
  1859 => x"1080d8f4",
  1860 => x"11555690",
  1861 => x"74708105",
  1862 => x"5681b72d",
  1863 => x"a07481b7",
  1864 => x"2d7681ff",
  1865 => x"06811658",
  1866 => x"5473802e",
  1867 => x"8a389c53",
  1868 => x"80d6b452",
  1869 => x"babe048b",
  1870 => x"5380d1c0",
  1871 => x"085280d8",
  1872 => x"f61651ba",
  1873 => x"f9047416",
  1874 => x"822bb8b9",
  1875 => x"0b80d090",
  1876 => x"120c5476",
  1877 => x"81ff0681",
  1878 => x"16585473",
  1879 => x"802e8a38",
  1880 => x"9c5380d6",
  1881 => x"b452baf0",
  1882 => x"048b5380",
  1883 => x"d1c00852",
  1884 => x"77753110",
  1885 => x"80d8f405",
  1886 => x"517655b7",
  1887 => x"bc2dbb96",
  1888 => x"04749029",
  1889 => x"75317010",
  1890 => x"80d8f405",
  1891 => x"515480d1",
  1892 => x"c0087481",
  1893 => x"b72d8119",
  1894 => x"59748b24",
  1895 => x"a338b9be",
  1896 => x"04749029",
  1897 => x"75317010",
  1898 => x"80d8f405",
  1899 => x"8c773157",
  1900 => x"51548074",
  1901 => x"81b72d9e",
  1902 => x"14ff1656",
  1903 => x"5474f338",
  1904 => x"02a4050d",
  1905 => x"0402fc05",
  1906 => x"0d80d1bc",
  1907 => x"081351b7",
  1908 => x"eb2d80d1",
  1909 => x"c008802e",
  1910 => x"893880d1",
  1911 => x"c00851a9",
  1912 => x"8a2d800b",
  1913 => x"80d1bc0c",
  1914 => x"b8f92d93",
  1915 => x"db2d0284",
  1916 => x"050d0402",
  1917 => x"fc050d72",
  1918 => x"5170fd2e",
  1919 => x"b03870fd",
  1920 => x"248a3870",
  1921 => x"fc2e80cc",
  1922 => x"38bcde04",
  1923 => x"70fe2eb7",
  1924 => x"3870ff2e",
  1925 => x"09810680",
  1926 => x"c53880d1",
  1927 => x"bc085170",
  1928 => x"802ebb38",
  1929 => x"ff1180d1",
  1930 => x"bc0cbcde",
  1931 => x"0480d1bc",
  1932 => x"08f40570",
  1933 => x"80d1bc0c",
  1934 => x"51708025",
  1935 => x"a138800b",
  1936 => x"80d1bc0c",
  1937 => x"bcde0480",
  1938 => x"d1bc0881",
  1939 => x"0580d1bc",
  1940 => x"0cbcde04",
  1941 => x"80d1bc08",
  1942 => x"8c0580d1",
  1943 => x"bc0cb8f9",
  1944 => x"2d93db2d",
  1945 => x"0284050d",
  1946 => x"0402fc05",
  1947 => x"0d800b80",
  1948 => x"d1bc0cb8",
  1949 => x"f92d92c9",
  1950 => x"2d80d1c0",
  1951 => x"0880d1ac",
  1952 => x"0c80d088",
  1953 => x"5195812d",
  1954 => x"0284050d",
  1955 => x"0402fc05",
  1956 => x"0d810b80",
  1957 => x"c8fc0c72",
  1958 => x"51bce92d",
  1959 => x"0284050d",
  1960 => x"0402fc05",
  1961 => x"0d800b80",
  1962 => x"c8fc0c72",
  1963 => x"51bce92d",
  1964 => x"0284050d",
  1965 => x"047180d8",
  1966 => x"f00c0400",
  1967 => x"00ffffff",
  1968 => x"ff00ffff",
  1969 => x"ffff00ff",
  1970 => x"ffffff00",
  1971 => x"4b455953",
  1972 => x"50312020",
  1973 => x"20202000",
  1974 => x"00000000",
  1975 => x"4b455953",
  1976 => x"50322020",
  1977 => x"20202000",
  1978 => x"00000000",
  1979 => x"3d3d2056",
  1980 => x"6964656f",
  1981 => x"70616320",
  1982 => x"666f7220",
  1983 => x"5a58444f",
  1984 => x"53203d3d",
  1985 => x"00000000",
  1986 => x"3d3d3d3d",
  1987 => x"3d3d3d3d",
  1988 => x"3d3d3d3d",
  1989 => x"3d3d3d3d",
  1990 => x"3d3d3d3d",
  1991 => x"3d3d3d3d",
  1992 => x"00000000",
  1993 => x"52657365",
  1994 => x"74000000",
  1995 => x"5363616e",
  1996 => x"6c696e65",
  1997 => x"73000000",
  1998 => x"53776170",
  1999 => x"206a6f79",
  2000 => x"73746963",
  2001 => x"6b730000",
  2002 => x"4a6f696e",
  2003 => x"206a6f79",
  2004 => x"73746963",
  2005 => x"6b730000",
  2006 => x"4c6f6164",
  2007 => x"20636174",
  2008 => x"72696467",
  2009 => x"6520524f",
  2010 => x"4d201000",
  2011 => x"4c6f6164",
  2012 => x"20564443",
  2013 => x"20666f6e",
  2014 => x"74201000",
  2015 => x"48656c70",
  2016 => x"00000000",
  2017 => x"45786974",
  2018 => x"00000000",
  2019 => x"54686520",
  2020 => x"766f6963",
  2021 => x"653a204f",
  2022 => x"66660000",
  2023 => x"54686520",
  2024 => x"766f6963",
  2025 => x"653a204f",
  2026 => x"6e000000",
  2027 => x"436f6c6f",
  2028 => x"72206d6f",
  2029 => x"64653a20",
  2030 => x"436f6c6f",
  2031 => x"72000000",
  2032 => x"436f6c6f",
  2033 => x"72206d6f",
  2034 => x"64653a20",
  2035 => x"4d6f6e6f",
  2036 => x"6368726f",
  2037 => x"6d650000",
  2038 => x"436f6c6f",
  2039 => x"72206d6f",
  2040 => x"64653a20",
  2041 => x"47726565",
  2042 => x"6e207068",
  2043 => x"6f737068",
  2044 => x"6f720000",
  2045 => x"436f6c6f",
  2046 => x"72206d6f",
  2047 => x"64653a20",
  2048 => x"416d6265",
  2049 => x"72206d6f",
  2050 => x"6e6f6368",
  2051 => x"726f6d65",
  2052 => x"00000000",
  2053 => x"4d6f6465",
  2054 => x"3a204f64",
  2055 => x"79737365",
  2056 => x"79322028",
  2057 => x"4e545343",
  2058 => x"29000000",
  2059 => x"4d6f6465",
  2060 => x"3a205669",
  2061 => x"64656f70",
  2062 => x"61632028",
  2063 => x"50414c29",
  2064 => x"00000000",
  2065 => x"3d3d2056",
  2066 => x"6964656f",
  2067 => x"70616320",
  2068 => x"666f7220",
  2069 => x"5a58554e",
  2070 => x"4f203d3d",
  2071 => x"00000000",
  2072 => x"5a58554e",
  2073 => x"4f3a2073",
  2074 => x"696e676c",
  2075 => x"65206a6f",
  2076 => x"79737469",
  2077 => x"636b0000",
  2078 => x"5a58554e",
  2079 => x"4f3a2032",
  2080 => x"206a6f79",
  2081 => x"73746963",
  2082 => x"6b207370",
  2083 => x"6c697474",
  2084 => x"65720000",
  2085 => x"5a58554e",
  2086 => x"4f3a2032",
  2087 => x"206a6f79",
  2088 => x"73746963",
  2089 => x"6b205647",
  2090 => x"41324d00",
  2091 => x"524f4d20",
  2092 => x"6c6f6164",
  2093 => x"696e6720",
  2094 => x"6661696c",
  2095 => x"65640000",
  2096 => x"4f4b0000",
  2097 => x"3d3d3d20",
  2098 => x"56696465",
  2099 => x"6f706163",
  2100 => x"20537065",
  2101 => x"6369616c",
  2102 => x"2048454c",
  2103 => x"50203d3d",
  2104 => x"3d000000",
  2105 => x"3d3d3d3d",
  2106 => x"3d3d3d3d",
  2107 => x"3d3d3d3d",
  2108 => x"3d3d3d3d",
  2109 => x"3d3d3d3d",
  2110 => x"3d3d3d3d",
  2111 => x"3d3d3d3d",
  2112 => x"3d3d0000",
  2113 => x"5363726f",
  2114 => x"6c6c204c",
  2115 => x"6f636b3a",
  2116 => x"20636861",
  2117 => x"6e676520",
  2118 => x"62657477",
  2119 => x"65656e00",
  2120 => x"52474220",
  2121 => x"616e6420",
  2122 => x"56474120",
  2123 => x"76696465",
  2124 => x"6f206d6f",
  2125 => x"64650000",
  2126 => x"46333a20",
  2127 => x"536f6674",
  2128 => x"20526573",
  2129 => x"65740000",
  2130 => x"4374726c",
  2131 => x"2b416c74",
  2132 => x"2b426163",
  2133 => x"6b737061",
  2134 => x"63653a20",
  2135 => x"48617264",
  2136 => x"20726573",
  2137 => x"65740000",
  2138 => x"45736320",
  2139 => x"6f72206a",
  2140 => x"6f797374",
  2141 => x"69636b20",
  2142 => x"62742e32",
  2143 => x"3a20746f",
  2144 => x"2073686f",
  2145 => x"77000000",
  2146 => x"6f722068",
  2147 => x"69646520",
  2148 => x"74686520",
  2149 => x"6f707469",
  2150 => x"6f6e7320",
  2151 => x"6d656e75",
  2152 => x"2e000000",
  2153 => x"57415344",
  2154 => x"202f2063",
  2155 => x"7572736f",
  2156 => x"72206b65",
  2157 => x"7973202f",
  2158 => x"206a6f79",
  2159 => x"73746963",
  2160 => x"6b000000",
  2161 => x"746f2073",
  2162 => x"656c6563",
  2163 => x"74206d65",
  2164 => x"6e75206f",
  2165 => x"7074696f",
  2166 => x"6e2e0000",
  2167 => x"456e7465",
  2168 => x"72202f20",
  2169 => x"46697265",
  2170 => x"20746f20",
  2171 => x"63686f6f",
  2172 => x"7365206f",
  2173 => x"7074696f",
  2174 => x"6e2e0000",
  2175 => x"496e206d",
  2176 => x"6f737420",
  2177 => x"67616d65",
  2178 => x"73207072",
  2179 => x"65737320",
  2180 => x"302d3920",
  2181 => x"61667465",
  2182 => x"72000000",
  2183 => x"6c6f6164",
  2184 => x"696e6720",
  2185 => x"6120524f",
  2186 => x"4d20746f",
  2187 => x"20706c61",
  2188 => x"79207468",
  2189 => x"65206761",
  2190 => x"6d650000",
  2191 => x"3d3d3d20",
  2192 => x"56696465",
  2193 => x"6f706163",
  2194 => x"20436f72",
  2195 => x"65204372",
  2196 => x"65646974",
  2197 => x"73203d3d",
  2198 => x"3d000000",
  2199 => x"3d3d3d3d",
  2200 => x"3d3d3d3d",
  2201 => x"3d3d3d3d",
  2202 => x"3d3d3d3d",
  2203 => x"3d3d3d3d",
  2204 => x"3d3d3d3d",
  2205 => x"3d3d3d3d",
  2206 => x"3d000000",
  2207 => x"5068696c",
  2208 => x"69707320",
  2209 => x"56696465",
  2210 => x"6f706163",
  2211 => x"202f204d",
  2212 => x"61676e61",
  2213 => x"766f7800",
  2214 => x"4f647973",
  2215 => x"73657932",
  2216 => x"20636f72",
  2217 => x"6520666f",
  2218 => x"72205a58",
  2219 => x"554e4f2c",
  2220 => x"205a5844",
  2221 => x"4f530000",
  2222 => x"616e6420",
  2223 => x"5a58444f",
  2224 => x"532b2062",
  2225 => x"6f617264",
  2226 => x"732e0000",
  2227 => x"4f726967",
  2228 => x"696e616c",
  2229 => x"20636f72",
  2230 => x"65206279",
  2231 => x"3a41726e",
  2232 => x"696d204c",
  2233 => x"61657567",
  2234 => x"65720000",
  2235 => x"506f7274",
  2236 => x"206d6164",
  2237 => x"65206279",
  2238 => x"3a20796f",
  2239 => x"6d626f70",
  2240 => x"72696d65",
  2241 => x"2c200000",
  2242 => x"2072616d",
  2243 => x"70613036",
  2244 => x"392c206e",
  2245 => x"6575726f",
  2246 => x"72756c65",
  2247 => x"7a2c2041",
  2248 => x"6e746f6e",
  2249 => x"696f0000",
  2250 => x"2053616e",
  2251 => x"6368657a",
  2252 => x"2c204176",
  2253 => x"6c697841",
  2254 => x"2c204d65",
  2255 => x"6a696173",
  2256 => x"33442c20",
  2257 => x"00000000",
  2258 => x"2057696c",
  2259 => x"636f3230",
  2260 => x"30392061",
  2261 => x"6e642042",
  2262 => x"656e6974",
  2263 => x"6f737300",
  2264 => x"53706563",
  2265 => x"69616c20",
  2266 => x"5468616e",
  2267 => x"6b732074",
  2268 => x"6f3a2052",
  2269 => x"656e6520",
  2270 => x"76616e20",
  2271 => x"00000000",
  2272 => x"2064656e",
  2273 => x"20456e64",
  2274 => x"656e2066",
  2275 => x"6f722068",
  2276 => x"69732069",
  2277 => x"6e666f20",
  2278 => x"6f6e2000",
  2279 => x"20766964",
  2280 => x"656f7061",
  2281 => x"632e6e6c",
  2282 => x"00000000",
  2283 => x"496e6974",
  2284 => x"69616c69",
  2285 => x"7a696e67",
  2286 => x"20534420",
  2287 => x"63617264",
  2288 => x"0a000000",
  2289 => x"16200000",
  2290 => x"14200000",
  2291 => x"15200000",
  2292 => x"53442069",
  2293 => x"6e69742e",
  2294 => x"2e2e0a00",
  2295 => x"53442063",
  2296 => x"61726420",
  2297 => x"72657365",
  2298 => x"74206661",
  2299 => x"696c6564",
  2300 => x"210a0000",
  2301 => x"53444843",
  2302 => x"20657272",
  2303 => x"6f72210a",
  2304 => x"00000000",
  2305 => x"57726974",
  2306 => x"65206661",
  2307 => x"696c6564",
  2308 => x"0a000000",
  2309 => x"52656164",
  2310 => x"20666169",
  2311 => x"6c65640a",
  2312 => x"00000000",
  2313 => x"43617264",
  2314 => x"20696e69",
  2315 => x"74206661",
  2316 => x"696c6564",
  2317 => x"0a000000",
  2318 => x"46415431",
  2319 => x"36202020",
  2320 => x"00000000",
  2321 => x"46415433",
  2322 => x"32202020",
  2323 => x"00000000",
  2324 => x"4e6f2070",
  2325 => x"61727469",
  2326 => x"74696f6e",
  2327 => x"20736967",
  2328 => x"0a000000",
  2329 => x"42616420",
  2330 => x"70617274",
  2331 => x"0a000000",
  2332 => x"4261636b",
  2333 => x"00000000",
  2334 => x"00000002",
  2335 => x"00000000",
  2336 => x"00000010",
  2337 => x"00000002",
  2338 => x"00001eec",
  2339 => x"000003ab",
  2340 => x"00000002",
  2341 => x"00001f08",
  2342 => x"000003ab",
  2343 => x"00000002",
  2344 => x"00001f24",
  2345 => x"0000037f",
  2346 => x"00000001",
  2347 => x"00001f2c",
  2348 => x"00000000",
  2349 => x"00000001",
  2350 => x"00001f38",
  2351 => x"00000001",
  2352 => x"00000001",
  2353 => x"00001f48",
  2354 => x"00000002",
  2355 => x"00000002",
  2356 => x"00001f58",
  2357 => x"00001ea1",
  2358 => x"00000002",
  2359 => x"00001f6c",
  2360 => x"00001e8d",
  2361 => x"00000003",
  2362 => x"00002544",
  2363 => x"00000002",
  2364 => x"00000003",
  2365 => x"00002534",
  2366 => x"00000004",
  2367 => x"00000003",
  2368 => x"0000252c",
  2369 => x"00000002",
  2370 => x"00000002",
  2371 => x"00001f7c",
  2372 => x"000003c6",
  2373 => x"00000002",
  2374 => x"00001f84",
  2375 => x"00000966",
  2376 => x"00000000",
  2377 => x"00000000",
  2378 => x"00000000",
  2379 => x"00001f8c",
  2380 => x"00001f9c",
  2381 => x"00001fac",
  2382 => x"00001fc0",
  2383 => x"00001fd8",
  2384 => x"00001ff4",
  2385 => x"00002014",
  2386 => x"0000202c",
  2387 => x"00000002",
  2388 => x"00002044",
  2389 => x"000003ab",
  2390 => x"00000002",
  2391 => x"00001f08",
  2392 => x"000003ab",
  2393 => x"00000002",
  2394 => x"00001f24",
  2395 => x"0000037f",
  2396 => x"00000001",
  2397 => x"00001f2c",
  2398 => x"00000000",
  2399 => x"00000001",
  2400 => x"00001f38",
  2401 => x"00000001",
  2402 => x"00000001",
  2403 => x"00001f48",
  2404 => x"00000002",
  2405 => x"00000002",
  2406 => x"00001f58",
  2407 => x"00001ea1",
  2408 => x"00000002",
  2409 => x"00001f6c",
  2410 => x"00001e8d",
  2411 => x"00000003",
  2412 => x"00002544",
  2413 => x"00000002",
  2414 => x"00000003",
  2415 => x"00002534",
  2416 => x"00000004",
  2417 => x"00000003",
  2418 => x"000025f4",
  2419 => x"00000003",
  2420 => x"00000002",
  2421 => x"00001f7c",
  2422 => x"000003c6",
  2423 => x"00000002",
  2424 => x"00001f84",
  2425 => x"00000966",
  2426 => x"00000000",
  2427 => x"00000000",
  2428 => x"00000000",
  2429 => x"00002060",
  2430 => x"00002078",
  2431 => x"00002094",
  2432 => x"00000004",
  2433 => x"000020ac",
  2434 => x"00002600",
  2435 => x"00000004",
  2436 => x"000020c0",
  2437 => x"000028e8",
  2438 => x"00000000",
  2439 => x"00000000",
  2440 => x"00000000",
  2441 => x"00000002",
  2442 => x"000020c4",
  2443 => x"000003aa",
  2444 => x"00000002",
  2445 => x"000020e4",
  2446 => x"000003aa",
  2447 => x"00000002",
  2448 => x"00002104",
  2449 => x"000003aa",
  2450 => x"00000002",
  2451 => x"00002120",
  2452 => x"000003aa",
  2453 => x"00000002",
  2454 => x"00002138",
  2455 => x"000003aa",
  2456 => x"00000002",
  2457 => x"00002148",
  2458 => x"000003aa",
  2459 => x"00000002",
  2460 => x"00002168",
  2461 => x"000003aa",
  2462 => x"00000002",
  2463 => x"00002188",
  2464 => x"000003aa",
  2465 => x"00000002",
  2466 => x"000021a4",
  2467 => x"000003aa",
  2468 => x"00000002",
  2469 => x"000021c4",
  2470 => x"000003aa",
  2471 => x"00000002",
  2472 => x"000021dc",
  2473 => x"000003aa",
  2474 => x"00000002",
  2475 => x"000021fc",
  2476 => x"000003aa",
  2477 => x"00000002",
  2478 => x"0000221c",
  2479 => x"000003aa",
  2480 => x"00000004",
  2481 => x"000020c0",
  2482 => x"000028e8",
  2483 => x"00000000",
  2484 => x"00000000",
  2485 => x"00000000",
  2486 => x"00000002",
  2487 => x"0000223c",
  2488 => x"000003aa",
  2489 => x"00000002",
  2490 => x"0000225c",
  2491 => x"000003aa",
  2492 => x"00000002",
  2493 => x"0000227c",
  2494 => x"000003aa",
  2495 => x"00000002",
  2496 => x"00002298",
  2497 => x"000003aa",
  2498 => x"00000002",
  2499 => x"000022b8",
  2500 => x"000003aa",
  2501 => x"00000002",
  2502 => x"000022cc",
  2503 => x"000003aa",
  2504 => x"00000002",
  2505 => x"000022ec",
  2506 => x"000003aa",
  2507 => x"00000002",
  2508 => x"00002308",
  2509 => x"000003aa",
  2510 => x"00000002",
  2511 => x"00002328",
  2512 => x"000003aa",
  2513 => x"00000002",
  2514 => x"00002348",
  2515 => x"000003aa",
  2516 => x"00000002",
  2517 => x"00002360",
  2518 => x"000003aa",
  2519 => x"00000002",
  2520 => x"00002380",
  2521 => x"000003aa",
  2522 => x"00000002",
  2523 => x"0000239c",
  2524 => x"000003aa",
  2525 => x"00000004",
  2526 => x"000020c0",
  2527 => x"000028e8",
  2528 => x"00000000",
  2529 => x"00000000",
  2530 => x"00000000",
  2531 => x"00000000",
  2532 => x"00000000",
  2533 => x"00000000",
  2534 => x"00000000",
  2535 => x"00000000",
  2536 => x"00000000",
  2537 => x"00000000",
  2538 => x"00000000",
  2539 => x"00000000",
  2540 => x"00000000",
  2541 => x"00000000",
  2542 => x"00000000",
  2543 => x"00000000",
  2544 => x"00000000",
  2545 => x"00000000",
  2546 => x"00000000",
  2547 => x"00000000",
  2548 => x"00000000",
  2549 => x"00000006",
  2550 => x"00000043",
  2551 => x"00000042",
  2552 => x"0000003b",
  2553 => x"0000004b",
  2554 => x"00000033",
  2555 => x"0000001d",
  2556 => x"0000001b",
  2557 => x"0000001c",
  2558 => x"00000023",
  2559 => x"0000002b",
  2560 => x"00000000",
  2561 => x"00000000",
  2562 => x"00000002",
  2563 => x"00002c74",
  2564 => x"00001c39",
  2565 => x"00000002",
  2566 => x"00002c92",
  2567 => x"00001c39",
  2568 => x"00000002",
  2569 => x"00002cb0",
  2570 => x"00001c39",
  2571 => x"00000002",
  2572 => x"00002cce",
  2573 => x"00001c39",
  2574 => x"00000002",
  2575 => x"00002cec",
  2576 => x"00001c39",
  2577 => x"00000002",
  2578 => x"00002d0a",
  2579 => x"00001c39",
  2580 => x"00000002",
  2581 => x"00002d28",
  2582 => x"00001c39",
  2583 => x"00000002",
  2584 => x"00002d46",
  2585 => x"00001c39",
  2586 => x"00000002",
  2587 => x"00002d64",
  2588 => x"00001c39",
  2589 => x"00000002",
  2590 => x"00002d82",
  2591 => x"00001c39",
  2592 => x"00000002",
  2593 => x"00002da0",
  2594 => x"00001c39",
  2595 => x"00000002",
  2596 => x"00002dbe",
  2597 => x"00001c39",
  2598 => x"00000002",
  2599 => x"00002ddc",
  2600 => x"00001c39",
  2601 => x"00000004",
  2602 => x"00002470",
  2603 => x"00000000",
  2604 => x"00000000",
  2605 => x"00000000",
  2606 => x"00001df3",
  2607 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

