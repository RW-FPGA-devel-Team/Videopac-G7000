library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity sp0256_al2_decoded is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of sp0256_al2_decoded is
	type rom is array(0 to  4047) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"18",X"01",X"00",X"19",X"01",X"00",X"1A",X"01",X"00",X"1B",X"01",X"00",X"1C",X"01",X"00",
		X"1D",X"0A",X"00",X"27",X"0A",X"00",X"31",X"01",X"00",X"32",X"03",X"00",X"35",X"03",X"00",X"38",
		X"03",X"00",X"3B",X"03",X"00",X"3E",X"01",X"00",X"3F",X"04",X"00",X"43",X"06",X"00",X"49",X"01",
		X"00",X"4A",X"04",X"00",X"4E",X"03",X"00",X"51",X"02",X"00",X"53",X"06",X"00",X"59",X"08",X"00",
		X"61",X"02",X"00",X"63",X"03",X"00",X"66",X"01",X"00",X"67",X"03",X"00",X"6A",X"06",X"00",X"70",
		X"01",X"00",X"71",X"03",X"00",X"74",X"02",X"00",X"76",X"01",X"00",X"77",X"01",X"00",X"78",X"03",
		X"00",X"7B",X"05",X"00",X"80",X"03",X"00",X"83",X"03",X"00",X"86",X"03",X"00",X"89",X"03",X"00",
		X"8C",X"04",X"00",X"90",X"02",X"00",X"92",X"03",X"00",X"95",X"01",X"00",X"96",X"03",X"00",X"99",
		X"04",X"00",X"9D",X"03",X"00",X"A0",X"04",X"00",X"A4",X"03",X"00",X"A7",X"03",X"00",X"AA",X"0D",
		X"00",X"B7",X"04",X"00",X"BB",X"04",X"00",X"BF",X"03",X"00",X"C2",X"09",X"00",X"CB",X"0A",X"00",
		X"D5",X"06",X"00",X"DB",X"02",X"00",X"DD",X"01",X"00",X"DE",X"06",X"00",X"E4",X"02",X"00",X"E6",
		X"09",X"00",X"EF",X"09",X"00",X"F8",X"08",X"01",X"00",X"03",X"01",X"03",X"03",X"01",X"06",X"03",
		X"01",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"07",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1F",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"01",X"40",X"5B",X"A0",X"60",X"B8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"00",X"C0",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"01",X"00",X"50",X"5B",X"A0",X"60",X"A8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"00",X"80",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"01",X"00",X"70",X"5B",X"A0",X"60",X"B0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"04",X"00",X"A0",X"5B",X"A0",X"60",X"B8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"02",X"01",X"C0",X"5B",X"A8",X"60",X"C0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"04",X"02",X"80",X"5B",X"A8",X"60",X"D0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"02",X"02",X"80",X"5B",X"A8",X"60",X"E0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"09",X"01",X"00",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"01",X"03",X"00",X"5B",X"B0",X"70",X"C8",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"01",X"02",X"80",X"5B",X"C8",X"70",X"B0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"03",X"00",X"5B",X"C8",X"70",X"B0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"02",X"80",X"5B",X"B0",X"70",X"C8",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"02",X"00",X"5B",X"C8",X"70",X"F8",X"70",X"B8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"02",X"80",X"5B",X"B0",X"70",X"D0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"03",X"03",X"80",X"5B",X"B0",X"70",X"F8",X"70",X"E0",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"01",X"03",X"00",X"5B",X"A8",X"70",X"E0",X"70",X"F8",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"03",X"02",X"80",X"5B",X"A0",X"70",X"E8",X"70",X"00",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"02",X"01",X"00",X"5B",X"A0",X"70",X"F0",X"70",X"00",X"60",X"18",X"50",X"3C",X"44",X"00",X"00",
		X"06",X"06",X"00",X"5B",X"00",X"50",X"28",X"50",X"40",X"50",X"F8",X"10",X"E8",X"58",X"AA",X"64",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"38",X"40",X"FC",X"04",X"CB",X"68",
		X"05",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"20",X"40",X"C5",X"62",
		X"0D",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"40",X"F4",X"2C",X"BF",X"3B",
		X"06",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"50",X"F8",X"44",X"CF",X"3A",
		X"04",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"18",X"42",X"FA",X"30",
		X"04",X"01",X"C0",X"5B",X"18",X"60",X"30",X"50",X"38",X"20",X"00",X"10",X"00",X"60",X"E6",X"38",
		X"04",X"01",X"40",X"5B",X"18",X"50",X"28",X"40",X"40",X"30",X"FC",X"68",X"E8",X"52",X"DD",X"16",
		X"07",X"00",X"38",X"5B",X"00",X"30",X"18",X"20",X"38",X"40",X"FC",X"60",X"E0",X"2A",X"A1",X"54",
		X"03",X"00",X"50",X"5B",X"08",X"30",X"20",X"30",X"20",X"10",X"FC",X"68",X"E8",X"1C",X"A2",X"50",
		X"09",X"00",X"60",X"5B",X"08",X"30",X"20",X"40",X"20",X"10",X"FC",X"68",X"E0",X"24",X"9B",X"5B",
		X"05",X"06",X"00",X"5B",X"00",X"50",X"10",X"20",X"30",X"50",X"E8",X"60",X"34",X"1E",X"A0",X"6E",
		X"05",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"28",X"1C",X"4E",X"F4",X"21",
		X"04",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"20",X"1C",X"44",X"EA",X"53",
		X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"1C",X"46",X"E7",X"5A",
		X"05",X"00",X"1C",X"5B",X"98",X"60",X"C0",X"60",X"E0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"03",X"00",X"50",X"5B",X"98",X"60",X"C0",X"60",X"E8",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"01",X"00",X"C0",X"5B",X"98",X"60",X"C0",X"60",X"E8",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"02",X"02",X"80",X"5B",X"A0",X"60",X"C0",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"01",X"01",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"02",X"02",X"00",X"5B",X"A0",X"60",X"B8",X"60",X"F0",X"50",X"0C",X"40",X"20",X"3C",X"32",X"2B",
		X"06",X"06",X"00",X"5B",X"F0",X"50",X"18",X"20",X"28",X"60",X"D0",X"60",X"28",X"18",X"A8",X"61",
		X"06",X"00",X"A0",X"5B",X"F0",X"50",X"C0",X"30",X"E0",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"05",X"00",X"C0",X"5B",X"F0",X"50",X"C0",X"30",X"E0",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"05",X"00",X"E0",X"5B",X"F0",X"50",X"E0",X"30",X"C8",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"04",X"01",X"40",X"5B",X"F0",X"50",X"E0",X"30",X"C8",X"20",X"00",X"10",X"20",X"44",X"00",X"00",
		X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"48",X"10",X"40",X"DF",X"3F",
		X"05",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"28",X"40",X"E8",X"3F",
		X"0C",X"00",X"A0",X"5B",X"08",X"30",X"18",X"30",X"38",X"40",X"EC",X"30",X"D4",X"2E",X"CB",X"20",
		X"03",X"02",X"80",X"5B",X"00",X"60",X"18",X"50",X"38",X"50",X"F4",X"08",X"DC",X"5E",X"A1",X"5C",
		X"03",X"06",X"00",X"5B",X"08",X"00",X"28",X"40",X"38",X"40",X"04",X"60",X"F0",X"66",X"A1",X"5A",
		X"03",X"06",X"00",X"5B",X"28",X"40",X"38",X"40",X"08",X"00",X"04",X"50",X"F4",X"62",X"A4",X"57",
		X"02",X"06",X"00",X"5B",X"08",X"10",X"28",X"50",X"38",X"40",X"04",X"48",X"F4",X"64",X"9A",X"62",
		X"03",X"06",X"00",X"5B",X"08",X"20",X"28",X"50",X"38",X"40",X"04",X"38",X"F8",X"60",X"96",X"66",
		X"04",X"04",X"00",X"5B",X"08",X"30",X"28",X"50",X"38",X"50",X"FC",X"20",X"F8",X"62",X"92",X"6E",
		X"04",X"01",X"40",X"5B",X"08",X"40",X"28",X"40",X"38",X"40",X"F8",X"60",X"F4",X"0C",X"90",X"71",
		X"03",X"03",X"00",X"5B",X"A0",X"70",X"E8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"01",X"03",X"00",X"5B",X"A0",X"70",X"F0",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"03",X"02",X"80",X"5B",X"A0",X"70",X"F0",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"01",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"F8",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"05",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"01",X"01",X"C0",X"5B",X"98",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"06",X"00",X"A0",X"5B",X"90",X"70",X"F8",X"60",X"00",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"02",X"00",X"70",X"5B",X"90",X"70",X"F8",X"60",X"F8",X"20",X"04",X"30",X"28",X"52",X"00",X"00",
		X"03",X"02",X"80",X"5B",X"90",X"70",X"E0",X"70",X"00",X"60",X"10",X"10",X"1C",X"56",X"3A",X"49",
		X"02",X"02",X"00",X"5B",X"98",X"70",X"E0",X"70",X"00",X"60",X"10",X"10",X"1C",X"56",X"3A",X"49",
		X"03",X"05",X"00",X"5B",X"98",X"60",X"F0",X"60",X"D8",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C",
		X"02",X"05",X"00",X"5B",X"D0",X"60",X"F0",X"60",X"A0",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C",
		X"02",X"04",X"00",X"5B",X"F0",X"60",X"C8",X"60",X"A0",X"60",X"1C",X"58",X"24",X"4E",X"39",X"2C",
		X"08",X"04",X"00",X"5B",X"20",X"50",X"18",X"20",X"40",X"30",X"F8",X"60",X"C0",X"60",X"B2",X"5A",
		X"03",X"05",X"00",X"5B",X"C8",X"60",X"B8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41",
		X"02",X"05",X"00",X"5B",X"C8",X"60",X"B8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41",
		X"02",X"05",X"00",X"5B",X"B8",X"60",X"C8",X"60",X"F8",X"60",X"14",X"28",X"1C",X"36",X"44",X"41",
		X"03",X"01",X"C0",X"5B",X"10",X"50",X"28",X"40",X"30",X"30",X"08",X"30",X"F0",X"64",X"8E",X"70",
		X"02",X"01",X"80",X"5B",X"10",X"50",X"28",X"50",X"38",X"30",X"04",X"28",X"F4",X"5E",X"8C",X"76",
		X"04",X"02",X"80",X"5B",X"08",X"30",X"28",X"40",X"30",X"20",X"08",X"40",X"F4",X"5C",X"90",X"70",
		X"01",X"04",X"00",X"5B",X"10",X"30",X"20",X"50",X"38",X"40",X"00",X"38",X"F0",X"5A",X"95",X"69",
		X"03",X"07",X"00",X"5B",X"20",X"40",X"28",X"40",X"18",X"10",X"00",X"48",X"F0",X"60",X"98",X"69",
		X"01",X"06",X"00",X"5B",X"18",X"30",X"28",X"40",X"20",X"10",X"00",X"48",X"F0",X"5E",X"9C",X"68",
		X"09",X"03",X"00",X"5B",X"F8",X"40",X"20",X"50",X"30",X"50",X"F0",X"20",X"DC",X"4C",X"AE",X"66",
		X"06",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"28",X"08",X"4E",X"EB",X"0C",
		X"06",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"38",X"0C",X"3E",X"F1",X"1A",
		X"02",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"E8",X"F2",X"03",X"3F",
		X"03",X"00",X"04",X"5B",X"F8",X"30",X"18",X"40",X"40",X"30",X"E4",X"20",X"18",X"04",X"88",X"76",
		X"01",X"03",X"00",X"5B",X"20",X"50",X"18",X"10",X"30",X"40",X"F8",X"78",X"E0",X"74",X"98",X"6C",
		X"14",X"00",X"28",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"30",X"10",X"24",X"E5",X"3B",
		X"08",X"02",X"80",X"5B",X"F8",X"70",X"20",X"50",X"28",X"50",X"C0",X"68",X"18",X"06",X"A4",X"5E",
		X"08",X"02",X"80",X"5B",X"F0",X"60",X"18",X"60",X"20",X"40",X"D8",X"60",X"20",X"0C",X"9D",X"61",
		X"04",X"03",X"00",X"5B",X"18",X"50",X"20",X"50",X"38",X"30",X"F0",X"60",X"D0",X"66",X"A6",X"53",
		X"07",X"02",X"00",X"5B",X"18",X"60",X"28",X"50",X"40",X"40",X"F0",X"60",X"C8",X"62",X"9D",X"61",
		X"08",X"01",X"C0",X"5B",X"B8",X"60",X"D0",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"05",X"01",X"00",X"5B",X"B0",X"60",X"C8",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"04",X"00",X"A0",X"5B",X"B0",X"60",X"C0",X"60",X"F8",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"04",X"00",X"80",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"07",X"00",X"28",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"50",X"0C",X"20",X"20",X"44",X"00",X"00",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"20",X"14",X"32",X"E7",X"23",
		X"03",X"06",X"00",X"5B",X"18",X"50",X"20",X"50",X"40",X"30",X"F8",X"60",X"E4",X"72",X"9D",X"5D",
		X"08",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"48",X"F4",X"42",X"EA",X"2A",
		X"03",X"01",X"40",X"5B",X"20",X"30",X"30",X"50",X"18",X"10",X"F8",X"68",X"E8",X"58",X"9C",X"68",
		X"06",X"00",X"20",X"5B",X"08",X"30",X"28",X"50",X"50",X"40",X"F0",X"48",X"C8",X"68",X"A8",X"47",
		X"06",X"00",X"E0",X"5B",X"10",X"40",X"28",X"40",X"50",X"50",X"F0",X"40",X"D0",X"1A",X"DE",X"3A",
		X"02",X"01",X"40",X"5B",X"F0",X"60",X"18",X"40",X"20",X"40",X"D0",X"68",X"2C",X"18",X"C7",X"25",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"30",X"FC",X"F0",X"FB",X"41",
		X"03",X"03",X"80",X"5B",X"10",X"40",X"20",X"60",X"38",X"30",X"F8",X"30",X"F4",X"5E",X"A1",X"5C",
		X"06",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1C",X"50",X"0C",X"0E",X"FB",X"5C",
		X"03",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"18",X"42",X"FA",X"56",
		X"12",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"18",X"18",X"4A",X"FC",X"5B",
		X"04",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"18",X"10",X"2E",X"F8",X"4C",
		X"07",X"01",X"40",X"5B",X"C0",X"30",X"E0",X"40",X"F8",X"60",X"14",X"58",X"24",X"48",X"00",X"00",
		X"0B",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"42",X"FE",X"3F",
		X"02",X"00",X"38",X"5B",X"08",X"40",X"20",X"30",X"38",X"30",X"DC",X"48",X"BC",X"58",X"A4",X"54",
		X"03",X"00",X"60",X"5B",X"D0",X"60",X"10",X"70",X"20",X"30",X"BC",X"60",X"1C",X"08",X"A1",X"5D",
		X"04",X"00",X"A0",X"5B",X"D0",X"50",X"10",X"60",X"18",X"50",X"BC",X"60",X"20",X"0E",X"A3",X"5C",
		X"11",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"38",X"04",X"28",X"E3",X"27",
		X"12",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"38",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"30",X"04",X"12",X"DE",X"56",
		X"02",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"28",X"F4",X"1E",X"DC",X"49",
		X"07",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"38",X"0C",X"62",X"E2",X"37",
		X"01",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"20",X"10",X"36",X"F9",X"44",
		X"09",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2C",X"28",X"0C",X"44",X"E7",X"1B",
		X"06",X"04",X"00",X"5B",X"20",X"50",X"40",X"60",X"58",X"50",X"00",X"58",X"DC",X"54",X"A7",X"4D",
		X"09",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"58",X"EC",X"00",X"21",X"30",
		X"04",X"05",X"00",X"5B",X"20",X"50",X"40",X"50",X"48",X"40",X"00",X"40",X"DC",X"60",X"B9",X"37",
		X"05",X"03",X"80",X"5B",X"D8",X"40",X"B8",X"40",X"F8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"03",X"02",X"00",X"5B",X"F0",X"40",X"B0",X"40",X"D8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"06",X"01",X"C0",X"5B",X"B0",X"40",X"F0",X"40",X"D8",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"08",X"01",X"40",X"5B",X"F0",X"40",X"B0",X"40",X"D0",X"40",X"04",X"58",X"2C",X"3C",X"55",X"5A",
		X"03",X"00",X"C0",X"5B",X"98",X"60",X"C8",X"60",X"08",X"40",X"18",X"30",X"28",X"44",X"2E",X"25",
		X"03",X"02",X"80",X"5B",X"A0",X"60",X"C8",X"60",X"08",X"40",X"18",X"30",X"28",X"44",X"2E",X"25",
		X"03",X"02",X"00",X"5B",X"A0",X"60",X"C0",X"60",X"00",X"40",X"18",X"30",X"28",X"44",X"2E",X"25",
		X"05",X"00",X"28",X"5B",X"F8",X"20",X"18",X"40",X"28",X"30",X"C0",X"38",X"10",X"F8",X"A0",X"5A",
		X"05",X"00",X"38",X"5B",X"08",X"30",X"20",X"60",X"38",X"40",X"FC",X"08",X"B0",X"50",X"9E",X"5F",
		X"06",X"00",X"50",X"5B",X"00",X"50",X"18",X"60",X"20",X"50",X"A8",X"70",X"14",X"02",X"93",X"72",
		X"03",X"02",X"80",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"02",X"80",X"5B",X"A0",X"60",X"E8",X"60",X"F8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"01",X"C0",X"5B",X"A0",X"60",X"E8",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"02",X"80",X"5B",X"A0",X"60",X"E0",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"03",X"00",X"5B",X"A8",X"60",X"E0",X"60",X"F0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"02",X"80",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"03",X"02",X"00",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"01",X"01",X"C0",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"03",X"00",X"E0",X"5B",X"A8",X"60",X"D0",X"60",X"E0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"01",X"00",X"80",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"02",X"00",X"C0",X"5B",X"A8",X"60",X"D0",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"01",X"00",X"70",X"5B",X"A8",X"60",X"D0",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"03",X"00",X"50",X"5B",X"A8",X"60",X"D8",X"60",X"E8",X"60",X"00",X"10",X"1C",X"52",X"42",X"59",
		X"06",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"FC",X"1C",X"D2",X"28",
		X"0B",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"38",X"04",X"18",X"B4",X"55",
		X"02",X"00",X"C0",X"5B",X"F8",X"40",X"30",X"70",X"20",X"20",X"C4",X"38",X"10",X"FC",X"A3",X"5D",
		X"02",X"01",X"40",X"5B",X"F8",X"60",X"28",X"50",X"28",X"50",X"B0",X"68",X"1C",X"06",X"A3",X"58",
		X"03",X"01",X"C0",X"5B",X"10",X"50",X"28",X"40",X"30",X"30",X"08",X"30",X"F0",X"64",X"8E",X"70",
		X"02",X"01",X"80",X"5B",X"10",X"50",X"28",X"50",X"38",X"30",X"04",X"28",X"F4",X"5E",X"8C",X"76",
		X"04",X"02",X"80",X"5B",X"08",X"30",X"28",X"40",X"30",X"20",X"08",X"40",X"F4",X"5C",X"90",X"70",
		X"01",X"04",X"00",X"5B",X"10",X"30",X"20",X"50",X"38",X"40",X"00",X"38",X"F0",X"5A",X"95",X"69",
		X"05",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"14",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"28",X"40",X"08",X"4E",X"E4",X"19",
		X"0D",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"34",X"50",X"10",X"66",X"F6",X"49",
		X"01",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"30",X"20",X"E4",X"60",X"CC",X"68",X"A5",X"5F",
		X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"28",X"10",X"E4",X"58",X"D0",X"60",X"A5",X"5F",
		X"01",X"02",X"80",X"5B",X"E0",X"60",X"18",X"40",X"20",X"40",X"D0",X"60",X"24",X"12",X"A8",X"5B",
		X"01",X"02",X"00",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"20",X"0A",X"A3",X"63",
		X"01",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D0",X"68",X"20",X"0A",X"A5",X"61",
		X"02",X"02",X"00",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"24",X"12",X"A2",X"69",
		X"01",X"01",X"40",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D4",X"68",X"1C",X"0A",X"A0",X"6E",
		X"02",X"00",X"E0",X"5B",X"18",X"60",X"20",X"20",X"20",X"10",X"E0",X"60",X"D4",X"68",X"A0",X"6E",
		X"01",X"01",X"00",X"5B",X"18",X"60",X"18",X"20",X"30",X"20",X"E4",X"60",X"D4",X"6A",X"A3",X"63",
		X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"30",X"20",X"E4",X"60",X"CC",X"68",X"A5",X"5F",
		X"02",X"02",X"80",X"5B",X"18",X"40",X"20",X"40",X"28",X"10",X"E4",X"58",X"D0",X"60",X"A5",X"5F",
		X"02",X"02",X"00",X"5B",X"E0",X"60",X"18",X"40",X"28",X"40",X"D0",X"60",X"24",X"10",X"A9",X"59",
		X"02",X"02",X"00",X"5B",X"E0",X"60",X"18",X"40",X"20",X"40",X"D0",X"60",X"24",X"12",X"A8",X"5B",
		X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"20",X"0A",X"A3",X"63",
		X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D0",X"68",X"20",X"0A",X"A5",X"61",
		X"02",X"01",X"C0",X"5B",X"E0",X"60",X"18",X"50",X"28",X"40",X"D0",X"60",X"24",X"12",X"A2",X"69",
		X"03",X"01",X"40",X"5B",X"E0",X"60",X"18",X"60",X"28",X"40",X"D4",X"68",X"1C",X"0A",X"A0",X"6E",
		X"03",X"00",X"C0",X"5B",X"18",X"60",X"20",X"20",X"20",X"10",X"E0",X"60",X"D4",X"68",X"A0",X"6E",
		X"03",X"00",X"E0",X"5B",X"18",X"60",X"18",X"20",X"30",X"20",X"E4",X"60",X"D4",X"6A",X"A3",X"63",
		X"03",X"02",X"80",X"5B",X"A8",X"60",X"C0",X"60",X"F8",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"03",X"02",X"00",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"01",X"01",X"C0",X"5B",X"A8",X"60",X"C0",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"05",X"00",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"01",X"00",X"C0",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"06",X"00",X"70",X"5B",X"A0",X"60",X"B8",X"60",X"00",X"60",X"40",X"60",X"24",X"60",X"00",X"00",
		X"11",X"00",X"A0",X"5B",X"08",X"30",X"18",X"30",X"38",X"40",X"EC",X"30",X"D4",X"2E",X"CB",X"20",
		X"03",X"02",X"80",X"5B",X"00",X"60",X"18",X"50",X"38",X"50",X"F4",X"08",X"DC",X"5E",X"A1",X"5C",
		X"0A",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"48",X"40",X"20",X"38",X"E3",X"29",
		X"04",X"00",X"A0",X"5B",X"00",X"30",X"18",X"20",X"38",X"40",X"FC",X"60",X"E0",X"2A",X"A1",X"54",
		X"02",X"00",X"C0",X"5B",X"08",X"30",X"20",X"30",X"20",X"10",X"FC",X"68",X"E8",X"1C",X"A2",X"50",
		X"02",X"00",X"C0",X"5B",X"08",X"30",X"20",X"40",X"20",X"10",X"FC",X"68",X"E0",X"24",X"9B",X"5B",
		X"03",X"06",X"00",X"5B",X"10",X"40",X"18",X"40",X"30",X"30",X"F8",X"68",X"DC",X"62",X"A8",X"50",
		X"01",X"06",X"00",X"5B",X"10",X"20",X"18",X"40",X"30",X"40",X"F8",X"68",X"D4",X"6E",X"AC",X"55",
		X"03",X"06",X"00",X"5B",X"20",X"50",X"18",X"10",X"30",X"40",X"F8",X"70",X"D0",X"6A",X"AC",X"58",
		X"0E",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"00",X"1E",X"C1",X"48",
		X"04",X"00",X"C0",X"5B",X"00",X"40",X"20",X"60",X"38",X"50",X"E8",X"18",X"E0",X"0A",X"C2",X"49",
		X"02",X"00",X"60",X"5B",X"A0",X"60",X"A8",X"60",X"F8",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"01",X"00",X"40",X"5B",X"A0",X"60",X"A8",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"03",X"00",X"50",X"5B",X"A0",X"60",X"A8",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"03",X"00",X"E0",X"5B",X"A0",X"60",X"B0",X"60",X"F0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"05",X"01",X"40",X"5B",X"A0",X"60",X"C0",X"60",X"E8",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"04",X"01",X"C0",X"5B",X"A8",X"60",X"C8",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"04",X"01",X"C0",X"5B",X"A8",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"01",X"00",X"E0",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"03",X"00",X"60",X"5B",X"A0",X"60",X"D0",X"60",X"E0",X"60",X"10",X"20",X"20",X"60",X"37",X"57",
		X"02",X"01",X"00",X"5B",X"18",X"60",X"28",X"40",X"10",X"00",X"F0",X"48",X"BC",X"64",X"AC",X"59",
		X"02",X"01",X"40",X"5B",X"10",X"60",X"20",X"40",X"18",X"10",X"F0",X"48",X"BC",X"62",X"AF",X"56",
		X"02",X"01",X"80",X"5B",X"10",X"50",X"20",X"30",X"20",X"10",X"EC",X"48",X"C0",X"5E",X"B0",X"56",
		X"02",X"01",X"40",X"5B",X"F0",X"50",X"10",X"60",X"20",X"50",X"C0",X"60",X"10",X"02",X"B6",X"51",
		X"02",X"01",X"40",X"5B",X"E8",X"60",X"18",X"60",X"28",X"50",X"C4",X"60",X"04",X"00",X"B8",X"4A",
		X"03",X"01",X"40",X"5B",X"18",X"60",X"10",X"00",X"20",X"30",X"E8",X"58",X"C8",X"62",X"B5",X"54",
		X"03",X"00",X"E0",X"5B",X"00",X"00",X"18",X"60",X"30",X"50",X"E4",X"60",X"CC",X"58",X"B5",X"56",
		X"03",X"00",X"C0",X"5B",X"00",X"00",X"18",X"60",X"28",X"40",X"E4",X"60",X"D0",X"5C",X"B2",X"59",
		X"03",X"00",X"80",X"5B",X"E8",X"60",X"10",X"60",X"20",X"20",X"CC",X"60",X"04",X"FC",X"B2",X"55",
		X"03",X"03",X"80",X"5B",X"90",X"70",X"F0",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"02",X"04",X"00",X"5B",X"90",X"70",X"F8",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"03",X"05",X"00",X"5B",X"90",X"70",X"F8",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"02",X"02",X"80",X"5B",X"90",X"70",X"F0",X"50",X"00",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"03",X"02",X"80",X"5B",X"98",X"70",X"E8",X"50",X"F8",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"04",X"01",X"80",X"5B",X"A0",X"70",X"E0",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"05",X"01",X"80",X"5B",X"A0",X"70",X"D8",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"05",X"01",X"40",X"5B",X"A0",X"70",X"D8",X"50",X"F0",X"30",X"04",X"18",X"28",X"4E",X"39",X"41",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"38",X"E0",X"40",X"E6",X"1C",
		X"02",X"01",X"80",X"5B",X"F8",X"40",X"18",X"60",X"38",X"50",X"F8",X"18",X"D8",X"5C",X"A1",X"70",
		X"05",X"03",X"00",X"5B",X"18",X"40",X"28",X"50",X"20",X"20",X"FC",X"68",X"C4",X"60",X"A3",X"64",
		X"03",X"01",X"80",X"5B",X"10",X"10",X"28",X"60",X"38",X"40",X"FC",X"60",X"C0",X"62",X"A3",X"60",
		X"07",X"01",X"00",X"5B",X"28",X"60",X"18",X"10",X"30",X"30",X"00",X"60",X"C0",X"60",X"A0",X"68",
		X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"30",X"FC",X"24",X"DE",X"43",
		X"02",X"05",X"00",X"5B",X"20",X"50",X"30",X"40",X"18",X"10",X"F8",X"68",X"E0",X"6E",X"99",X"6C");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
