-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb8",
     9 => x"c0080b0b",
    10 => x"0bb8c408",
    11 => x"0b0b0bb8",
    12 => x"c8080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b8c80c0b",
    16 => x"0b0bb8c4",
    17 => x"0c0b0b0b",
    18 => x"b8c00c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafa4",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b8c07080",
    57 => x"c2f0278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e604",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb8d00c",
    65 => x"9f0bb8d4",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b8d408ff",
    69 => x"05b8d40c",
    70 => x"b8d40880",
    71 => x"25eb38b8",
    72 => x"d008ff05",
    73 => x"b8d00cb8",
    74 => x"d0088025",
    75 => x"d738800b",
    76 => x"b8d40c80",
    77 => x"0bb8d00c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb8d008",
    97 => x"258f3882",
    98 => x"bd2db8d0",
    99 => x"08ff05b8",
   100 => x"d00c82ff",
   101 => x"04b8d008",
   102 => x"b8d40853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b8d008a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b8d4",
   111 => x"088105b8",
   112 => x"d40cb8d4",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb8d40c",
   116 => x"b8d00881",
   117 => x"05b8d00c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b8",
   122 => x"d4088105",
   123 => x"b8d40cb8",
   124 => x"d408a02e",
   125 => x"0981068e",
   126 => x"38800bb8",
   127 => x"d40cb8d0",
   128 => x"088105b8",
   129 => x"d00c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb8d8",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb8d80c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b8",
   169 => x"d8088407",
   170 => x"b8d80c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb4c0",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b8d80852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b8c00c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c8dc12d",
   216 => x"0284050d",
   217 => x"0402fc05",
   218 => x"0dec5192",
   219 => x"710c86a4",
   220 => x"2d82710c",
   221 => x"0284050d",
   222 => x"0402d005",
   223 => x"0d7d5480",
   224 => x"5ba40bec",
   225 => x"0c7352b8",
   226 => x"dc51a6e0",
   227 => x"2db8c008",
   228 => x"7b2e81ab",
   229 => x"38b8e008",
   230 => x"70f80c89",
   231 => x"1580f52d",
   232 => x"8a1680f5",
   233 => x"2d718280",
   234 => x"29058817",
   235 => x"80f52d70",
   236 => x"84808029",
   237 => x"12f40c7e",
   238 => x"ff155c5e",
   239 => x"57555658",
   240 => x"767b2e8b",
   241 => x"38811a77",
   242 => x"812a585a",
   243 => x"76f738f7",
   244 => x"1a5a815b",
   245 => x"80782580",
   246 => x"e6387952",
   247 => x"7651848b",
   248 => x"2db9a852",
   249 => x"b8dc51a9",
   250 => x"962db8c0",
   251 => x"08802eb8",
   252 => x"38b9a85c",
   253 => x"83fc597b",
   254 => x"7084055d",
   255 => x"087081ff",
   256 => x"0671882a",
   257 => x"7081ff06",
   258 => x"73902a70",
   259 => x"81ff0675",
   260 => x"982ae80c",
   261 => x"e80c58e8",
   262 => x"0c57e80c",
   263 => x"fc1a5a53",
   264 => x"788025d3",
   265 => x"3888af04",
   266 => x"b8c0085b",
   267 => x"848058b8",
   268 => x"dc51a8e9",
   269 => x"2dfc8018",
   270 => x"81185858",
   271 => x"87d40486",
   272 => x"b72d800b",
   273 => x"ec0c7a80",
   274 => x"2e8d38b4",
   275 => x"c4518fbe",
   276 => x"2d8dc12d",
   277 => x"88dd04b6",
   278 => x"90518fbe",
   279 => x"2d7ab8c0",
   280 => x"0c02b005",
   281 => x"0d0402ec",
   282 => x"050d850b",
   283 => x"ec0c8da2",
   284 => x"2d8a8c2d",
   285 => x"81f82d9d",
   286 => x"fd2db8c0",
   287 => x"08802e80",
   288 => x"f63886f9",
   289 => x"51af9d2d",
   290 => x"b4c4518f",
   291 => x"be2d8dc1",
   292 => x"2d8a982d",
   293 => x"8fce2db4",
   294 => x"f00b80f5",
   295 => x"2d70892b",
   296 => x"9c8006b4",
   297 => x"fc0b80f5",
   298 => x"2d70872b",
   299 => x"818006b5",
   300 => x"880b80f5",
   301 => x"2d701082",
   302 => x"06747307",
   303 => x"07b5940b",
   304 => x"80f52d70",
   305 => x"8c2b81e0",
   306 => x"8006b5a0",
   307 => x"0b80f52d",
   308 => x"708f2b82",
   309 => x"80800674",
   310 => x"730707fc",
   311 => x"0c545456",
   312 => x"54525757",
   313 => x"54528652",
   314 => x"b8c00885",
   315 => x"38b8c008",
   316 => x"5271ec0c",
   317 => x"89910480",
   318 => x"0bb8c00c",
   319 => x"0294050d",
   320 => x"0471980c",
   321 => x"04ffb008",
   322 => x"b8c00c04",
   323 => x"810bffb0",
   324 => x"0c04800b",
   325 => x"ffb00c04",
   326 => x"02f4050d",
   327 => x"8b9a04b8",
   328 => x"c00881f0",
   329 => x"2e098106",
   330 => x"8938810b",
   331 => x"b6f40c8b",
   332 => x"9a04b8c0",
   333 => x"0881e02e",
   334 => x"09810689",
   335 => x"38810bb6",
   336 => x"f80c8b9a",
   337 => x"04b8c008",
   338 => x"52b6f808",
   339 => x"802e8838",
   340 => x"b8c00881",
   341 => x"80055271",
   342 => x"842c728f",
   343 => x"065353b6",
   344 => x"f408802e",
   345 => x"99387284",
   346 => x"29b6b405",
   347 => x"72138171",
   348 => x"2b700973",
   349 => x"0806730c",
   350 => x"5153538b",
   351 => x"90047284",
   352 => x"29b6b405",
   353 => x"72138371",
   354 => x"2b720807",
   355 => x"720c5353",
   356 => x"800bb6f8",
   357 => x"0c800bb6",
   358 => x"f40cb8e8",
   359 => x"518c9b2d",
   360 => x"b8c008ff",
   361 => x"24fef838",
   362 => x"800bb8c0",
   363 => x"0c028c05",
   364 => x"0d0402f8",
   365 => x"050db6b4",
   366 => x"528f5180",
   367 => x"72708405",
   368 => x"540cff11",
   369 => x"51708025",
   370 => x"f2380288",
   371 => x"050d0402",
   372 => x"f0050d75",
   373 => x"518a922d",
   374 => x"70822cfc",
   375 => x"06b6b411",
   376 => x"72109e06",
   377 => x"71087072",
   378 => x"2a708306",
   379 => x"82742b70",
   380 => x"09740676",
   381 => x"0c545156",
   382 => x"57535153",
   383 => x"8a8c2d71",
   384 => x"b8c00c02",
   385 => x"90050d04",
   386 => x"02fc050d",
   387 => x"72518071",
   388 => x"0c800b84",
   389 => x"120c0284",
   390 => x"050d0402",
   391 => x"f0050d75",
   392 => x"70088412",
   393 => x"08535353",
   394 => x"ff547171",
   395 => x"2ea8388a",
   396 => x"922d8413",
   397 => x"08708429",
   398 => x"14881170",
   399 => x"087081ff",
   400 => x"06841808",
   401 => x"81118706",
   402 => x"841a0c53",
   403 => x"51555151",
   404 => x"518a8c2d",
   405 => x"715473b8",
   406 => x"c00c0290",
   407 => x"050d0402",
   408 => x"f8050d8a",
   409 => x"922de008",
   410 => x"708b2a70",
   411 => x"81065152",
   412 => x"5270802e",
   413 => x"9d38b8e8",
   414 => x"08708429",
   415 => x"b8f00573",
   416 => x"81ff0671",
   417 => x"0c5151b8",
   418 => x"e8088111",
   419 => x"8706b8e8",
   420 => x"0c51800b",
   421 => x"b9900c8a",
   422 => x"852d8a8c",
   423 => x"2d028805",
   424 => x"0d0402fc",
   425 => x"050db8e8",
   426 => x"518c882d",
   427 => x"8bb22d8c",
   428 => x"df518a81",
   429 => x"2d028405",
   430 => x"0d04b994",
   431 => x"08b8c00c",
   432 => x"0402fc05",
   433 => x"0d8dcb04",
   434 => x"8a982d80",
   435 => x"f6518bcf",
   436 => x"2db8c008",
   437 => x"f33880da",
   438 => x"518bcf2d",
   439 => x"b8c008e8",
   440 => x"38b8c008",
   441 => x"b7800cb8",
   442 => x"c0085184",
   443 => x"f02d0284",
   444 => x"050d0402",
   445 => x"ec050d76",
   446 => x"54805287",
   447 => x"0b881580",
   448 => x"f52d5653",
   449 => x"74722483",
   450 => x"38a05372",
   451 => x"5182f92d",
   452 => x"81128b15",
   453 => x"80f52d54",
   454 => x"52727225",
   455 => x"de380294",
   456 => x"050d0402",
   457 => x"f0050db9",
   458 => x"94085481",
   459 => x"f82d800b",
   460 => x"b9980c73",
   461 => x"08802e81",
   462 => x"8038820b",
   463 => x"b8d40cb9",
   464 => x"98088f06",
   465 => x"b8d00c73",
   466 => x"08527183",
   467 => x"2e963871",
   468 => x"83268938",
   469 => x"71812eaf",
   470 => x"388fa404",
   471 => x"71852e9f",
   472 => x"388fa404",
   473 => x"881480f5",
   474 => x"2d841508",
   475 => x"b38c5354",
   476 => x"5285fe2d",
   477 => x"71842913",
   478 => x"70085252",
   479 => x"8fa80473",
   480 => x"518df32d",
   481 => x"8fa404b6",
   482 => x"fc088815",
   483 => x"082c7081",
   484 => x"06515271",
   485 => x"802e8738",
   486 => x"b390518f",
   487 => x"a104b394",
   488 => x"5185fe2d",
   489 => x"84140851",
   490 => x"85fe2db9",
   491 => x"98088105",
   492 => x"b9980c8c",
   493 => x"14548eb3",
   494 => x"04029005",
   495 => x"0d0471b9",
   496 => x"940c8ea3",
   497 => x"2db99808",
   498 => x"ff05b99c",
   499 => x"0c0402e8",
   500 => x"050db994",
   501 => x"08b9a008",
   502 => x"57558751",
   503 => x"8bcf2db8",
   504 => x"c008812a",
   505 => x"70810651",
   506 => x"5271802e",
   507 => x"a0388ff4",
   508 => x"048a982d",
   509 => x"87518bcf",
   510 => x"2db8c008",
   511 => x"f438b780",
   512 => x"08813270",
   513 => x"b7800c70",
   514 => x"525284f0",
   515 => x"2d80fe51",
   516 => x"8bcf2db8",
   517 => x"c008802e",
   518 => x"a638b780",
   519 => x"08802e91",
   520 => x"38800bb7",
   521 => x"800c8051",
   522 => x"84f02d90",
   523 => x"b1048a98",
   524 => x"2d80fe51",
   525 => x"8bcf2db8",
   526 => x"c008f338",
   527 => x"86e52db7",
   528 => x"80089038",
   529 => x"81fd518b",
   530 => x"cf2d81fa",
   531 => x"518bcf2d",
   532 => x"96840481",
   533 => x"f5518bcf",
   534 => x"2db8c008",
   535 => x"812a7081",
   536 => x"06515271",
   537 => x"802eaf38",
   538 => x"b99c0852",
   539 => x"71802e89",
   540 => x"38ff12b9",
   541 => x"9c0c9196",
   542 => x"04b99808",
   543 => x"10b99808",
   544 => x"05708429",
   545 => x"16515288",
   546 => x"1208802e",
   547 => x"8938ff51",
   548 => x"88120852",
   549 => x"712d81f2",
   550 => x"518bcf2d",
   551 => x"b8c00881",
   552 => x"2a708106",
   553 => x"51527180",
   554 => x"2eb138b9",
   555 => x"9808ff11",
   556 => x"b99c0856",
   557 => x"53537372",
   558 => x"25893881",
   559 => x"14b99c0c",
   560 => x"91db0472",
   561 => x"10137084",
   562 => x"29165152",
   563 => x"88120880",
   564 => x"2e8938fe",
   565 => x"51881208",
   566 => x"52712d81",
   567 => x"fd518bcf",
   568 => x"2db8c008",
   569 => x"812a7081",
   570 => x"06515271",
   571 => x"802ead38",
   572 => x"b99c0880",
   573 => x"2e893880",
   574 => x"0bb99c0c",
   575 => x"929c04b9",
   576 => x"980810b9",
   577 => x"98080570",
   578 => x"84291651",
   579 => x"52881208",
   580 => x"802e8938",
   581 => x"fd518812",
   582 => x"0852712d",
   583 => x"81fa518b",
   584 => x"cf2db8c0",
   585 => x"08812a70",
   586 => x"81065152",
   587 => x"71802eae",
   588 => x"38b99808",
   589 => x"ff115452",
   590 => x"b99c0873",
   591 => x"25883872",
   592 => x"b99c0c92",
   593 => x"de047110",
   594 => x"12708429",
   595 => x"16515288",
   596 => x"1208802e",
   597 => x"8938fc51",
   598 => x"88120852",
   599 => x"712db99c",
   600 => x"08705354",
   601 => x"73802e8a",
   602 => x"388c15ff",
   603 => x"15555592",
   604 => x"e404820b",
   605 => x"b8d40c71",
   606 => x"8f06b8d0",
   607 => x"0c81eb51",
   608 => x"8bcf2db8",
   609 => x"c008812a",
   610 => x"70810651",
   611 => x"5271802e",
   612 => x"ad387408",
   613 => x"852e0981",
   614 => x"06a43888",
   615 => x"1580f52d",
   616 => x"ff055271",
   617 => x"881681b7",
   618 => x"2d71982b",
   619 => x"52718025",
   620 => x"8838800b",
   621 => x"881681b7",
   622 => x"2d74518d",
   623 => x"f32d81f4",
   624 => x"518bcf2d",
   625 => x"b8c00881",
   626 => x"2a708106",
   627 => x"51527180",
   628 => x"2eb33874",
   629 => x"08852e09",
   630 => x"8106aa38",
   631 => x"881580f5",
   632 => x"2d810552",
   633 => x"71881681",
   634 => x"b72d7181",
   635 => x"ff068b16",
   636 => x"80f52d54",
   637 => x"52727227",
   638 => x"87387288",
   639 => x"1681b72d",
   640 => x"74518df3",
   641 => x"2d80da51",
   642 => x"8bcf2db8",
   643 => x"c008812a",
   644 => x"70810651",
   645 => x"5271802e",
   646 => x"81a638b9",
   647 => x"9408b99c",
   648 => x"08555373",
   649 => x"802e8a38",
   650 => x"8c13ff15",
   651 => x"555394a3",
   652 => x"04720852",
   653 => x"71822ea6",
   654 => x"38718226",
   655 => x"89387181",
   656 => x"2ea93895",
   657 => x"c0047183",
   658 => x"2eb13871",
   659 => x"842e0981",
   660 => x"0680ed38",
   661 => x"88130851",
   662 => x"8fbe2d95",
   663 => x"c004b99c",
   664 => x"08518813",
   665 => x"0852712d",
   666 => x"95c00481",
   667 => x"0b881408",
   668 => x"2bb6fc08",
   669 => x"32b6fc0c",
   670 => x"95960488",
   671 => x"1380f52d",
   672 => x"81058b14",
   673 => x"80f52d53",
   674 => x"54717424",
   675 => x"83388054",
   676 => x"73881481",
   677 => x"b72d8ea3",
   678 => x"2d95c004",
   679 => x"7508802e",
   680 => x"a2387508",
   681 => x"518bcf2d",
   682 => x"b8c00881",
   683 => x"06527180",
   684 => x"2e8b38b9",
   685 => x"9c085184",
   686 => x"16085271",
   687 => x"2d881656",
   688 => x"75da3880",
   689 => x"54800bb8",
   690 => x"d40c738f",
   691 => x"06b8d00c",
   692 => x"a05273b9",
   693 => x"9c082e09",
   694 => x"81069838",
   695 => x"b99808ff",
   696 => x"05743270",
   697 => x"09810570",
   698 => x"72079f2a",
   699 => x"91713151",
   700 => x"51535371",
   701 => x"5182f92d",
   702 => x"8114548e",
   703 => x"7425c638",
   704 => x"b7800852",
   705 => x"71b8c00c",
   706 => x"0298050d",
   707 => x"0402f405",
   708 => x"0dd45281",
   709 => x"ff720c71",
   710 => x"085381ff",
   711 => x"720c7288",
   712 => x"2b83fe80",
   713 => x"06720870",
   714 => x"81ff0651",
   715 => x"525381ff",
   716 => x"720c7271",
   717 => x"07882b72",
   718 => x"087081ff",
   719 => x"06515253",
   720 => x"81ff720c",
   721 => x"72710788",
   722 => x"2b720870",
   723 => x"81ff0672",
   724 => x"07b8c00c",
   725 => x"5253028c",
   726 => x"050d0402",
   727 => x"f4050d74",
   728 => x"767181ff",
   729 => x"06d40c53",
   730 => x"53b9a408",
   731 => x"85387189",
   732 => x"2b527198",
   733 => x"2ad40c71",
   734 => x"902a7081",
   735 => x"ff06d40c",
   736 => x"5171882a",
   737 => x"7081ff06",
   738 => x"d40c5171",
   739 => x"81ff06d4",
   740 => x"0c72902a",
   741 => x"7081ff06",
   742 => x"d40c51d4",
   743 => x"087081ff",
   744 => x"06515182",
   745 => x"b8bf5270",
   746 => x"81ff2e09",
   747 => x"81069438",
   748 => x"81ff0bd4",
   749 => x"0cd40870",
   750 => x"81ff06ff",
   751 => x"14545151",
   752 => x"71e53870",
   753 => x"b8c00c02",
   754 => x"8c050d04",
   755 => x"02fc050d",
   756 => x"81c75181",
   757 => x"ff0bd40c",
   758 => x"ff115170",
   759 => x"8025f438",
   760 => x"0284050d",
   761 => x"0402f405",
   762 => x"0d81ff0b",
   763 => x"d40c9353",
   764 => x"805287fc",
   765 => x"80c15196",
   766 => x"db2db8c0",
   767 => x"088b3881",
   768 => x"ff0bd40c",
   769 => x"81539892",
   770 => x"0497cc2d",
   771 => x"ff135372",
   772 => x"df3872b8",
   773 => x"c00c028c",
   774 => x"050d0402",
   775 => x"ec050d81",
   776 => x"0bb9a40c",
   777 => x"8454d008",
   778 => x"708f2a70",
   779 => x"81065151",
   780 => x"5372f338",
   781 => x"72d00c97",
   782 => x"cc2db398",
   783 => x"5185fe2d",
   784 => x"d008708f",
   785 => x"2a708106",
   786 => x"51515372",
   787 => x"f338810b",
   788 => x"d00cb153",
   789 => x"805284d4",
   790 => x"80c05196",
   791 => x"db2db8c0",
   792 => x"08812e93",
   793 => x"3872822e",
   794 => x"bd38ff13",
   795 => x"5372e538",
   796 => x"ff145473",
   797 => x"ffb03897",
   798 => x"cc2d83aa",
   799 => x"52849c80",
   800 => x"c85196db",
   801 => x"2db8c008",
   802 => x"812e0981",
   803 => x"06923896",
   804 => x"8d2db8c0",
   805 => x"0883ffff",
   806 => x"06537283",
   807 => x"aa2e9d38",
   808 => x"97e52d99",
   809 => x"b704b3a4",
   810 => x"5185fe2d",
   811 => x"80539b85",
   812 => x"04b3bc51",
   813 => x"85fe2d80",
   814 => x"549ad704",
   815 => x"81ff0bd4",
   816 => x"0cb15497",
   817 => x"cc2d8fcf",
   818 => x"53805287",
   819 => x"fc80f751",
   820 => x"96db2db8",
   821 => x"c00855b8",
   822 => x"c008812e",
   823 => x"0981069b",
   824 => x"3881ff0b",
   825 => x"d40c820a",
   826 => x"52849c80",
   827 => x"e95196db",
   828 => x"2db8c008",
   829 => x"802e8d38",
   830 => x"97cc2dff",
   831 => x"135372c9",
   832 => x"389aca04",
   833 => x"81ff0bd4",
   834 => x"0cb8c008",
   835 => x"5287fc80",
   836 => x"fa5196db",
   837 => x"2db8c008",
   838 => x"b13881ff",
   839 => x"0bd40cd4",
   840 => x"085381ff",
   841 => x"0bd40c81",
   842 => x"ff0bd40c",
   843 => x"81ff0bd4",
   844 => x"0c81ff0b",
   845 => x"d40c7286",
   846 => x"2a708106",
   847 => x"76565153",
   848 => x"729538b8",
   849 => x"c008549a",
   850 => x"d7047382",
   851 => x"2efee238",
   852 => x"ff145473",
   853 => x"feed3873",
   854 => x"b9a40c73",
   855 => x"8b388152",
   856 => x"87fc80d0",
   857 => x"5196db2d",
   858 => x"81ff0bd4",
   859 => x"0cd00870",
   860 => x"8f2a7081",
   861 => x"06515153",
   862 => x"72f33872",
   863 => x"d00c81ff",
   864 => x"0bd40c81",
   865 => x"5372b8c0",
   866 => x"0c029405",
   867 => x"0d0402e8",
   868 => x"050d7855",
   869 => x"805681ff",
   870 => x"0bd40cd0",
   871 => x"08708f2a",
   872 => x"70810651",
   873 => x"515372f3",
   874 => x"3882810b",
   875 => x"d00c81ff",
   876 => x"0bd40c77",
   877 => x"5287fc80",
   878 => x"d15196db",
   879 => x"2d80dbc6",
   880 => x"df54b8c0",
   881 => x"08802e8a",
   882 => x"38b3dc51",
   883 => x"85fe2d9c",
   884 => x"a50481ff",
   885 => x"0bd40cd4",
   886 => x"087081ff",
   887 => x"06515372",
   888 => x"81fe2e09",
   889 => x"81069d38",
   890 => x"80ff5396",
   891 => x"8d2db8c0",
   892 => x"08757084",
   893 => x"05570cff",
   894 => x"13537280",
   895 => x"25ed3881",
   896 => x"569c8a04",
   897 => x"ff145473",
   898 => x"c93881ff",
   899 => x"0bd40c81",
   900 => x"ff0bd40c",
   901 => x"d008708f",
   902 => x"2a708106",
   903 => x"51515372",
   904 => x"f33872d0",
   905 => x"0c75b8c0",
   906 => x"0c029805",
   907 => x"0d0402e8",
   908 => x"050d7779",
   909 => x"7b585555",
   910 => x"80537276",
   911 => x"25a33874",
   912 => x"70810556",
   913 => x"80f52d74",
   914 => x"70810556",
   915 => x"80f52d52",
   916 => x"5271712e",
   917 => x"86388151",
   918 => x"9ce30481",
   919 => x"13539cba",
   920 => x"04805170",
   921 => x"b8c00c02",
   922 => x"98050d04",
   923 => x"02ec050d",
   924 => x"76557480",
   925 => x"2ebb389a",
   926 => x"1580e02d",
   927 => x"51a9ec2d",
   928 => x"b8c008b8",
   929 => x"c008bfd8",
   930 => x"0cb8c008",
   931 => x"5454bfb4",
   932 => x"08802e99",
   933 => x"38941580",
   934 => x"e02d51a9",
   935 => x"ec2db8c0",
   936 => x"08902b83",
   937 => x"fff00a06",
   938 => x"70750751",
   939 => x"5372bfd8",
   940 => x"0cbfd808",
   941 => x"5372802e",
   942 => x"9938bfac",
   943 => x"08fe1471",
   944 => x"29bfc008",
   945 => x"05bfdc0c",
   946 => x"70842bbf",
   947 => x"b80c549d",
   948 => x"f804bfc4",
   949 => x"08bfd80c",
   950 => x"bfc808bf",
   951 => x"dc0cbfb4",
   952 => x"08802e8a",
   953 => x"38bfac08",
   954 => x"842b539d",
   955 => x"f404bfcc",
   956 => x"08842b53",
   957 => x"72bfb80c",
   958 => x"0294050d",
   959 => x"0402d805",
   960 => x"0d800bbf",
   961 => x"b40c8454",
   962 => x"989b2db8",
   963 => x"c008802e",
   964 => x"9538b9a8",
   965 => x"5280519b",
   966 => x"8e2db8c0",
   967 => x"08802e86",
   968 => x"38fe549e",
   969 => x"ae04ff14",
   970 => x"54738024",
   971 => x"db38738c",
   972 => x"38b3ec51",
   973 => x"85fe2d73",
   974 => x"55a3b704",
   975 => x"8056810b",
   976 => x"bfe00c88",
   977 => x"53b48052",
   978 => x"b9de519c",
   979 => x"ae2db8c0",
   980 => x"08762e09",
   981 => x"81068738",
   982 => x"b8c008bf",
   983 => x"e00c8853",
   984 => x"b48c52b9",
   985 => x"fa519cae",
   986 => x"2db8c008",
   987 => x"8738b8c0",
   988 => x"08bfe00c",
   989 => x"bfe00880",
   990 => x"2e80f638",
   991 => x"bcee0b80",
   992 => x"f52dbcef",
   993 => x"0b80f52d",
   994 => x"71982b71",
   995 => x"902b07bc",
   996 => x"f00b80f5",
   997 => x"2d70882b",
   998 => x"7207bcf1",
   999 => x"0b80f52d",
  1000 => x"7107bda6",
  1001 => x"0b80f52d",
  1002 => x"bda70b80",
  1003 => x"f52d7188",
  1004 => x"2b07535f",
  1005 => x"54525a56",
  1006 => x"57557381",
  1007 => x"abaa2e09",
  1008 => x"81068d38",
  1009 => x"7551a9bc",
  1010 => x"2db8c008",
  1011 => x"569fdd04",
  1012 => x"7382d4d5",
  1013 => x"2e8738b4",
  1014 => x"9851a09e",
  1015 => x"04b9a852",
  1016 => x"75519b8e",
  1017 => x"2db8c008",
  1018 => x"55b8c008",
  1019 => x"802e83c7",
  1020 => x"388853b4",
  1021 => x"8c52b9fa",
  1022 => x"519cae2d",
  1023 => x"b8c00889",
  1024 => x"38810bbf",
  1025 => x"b40ca0a4",
  1026 => x"048853b4",
  1027 => x"8052b9de",
  1028 => x"519cae2d",
  1029 => x"b8c00880",
  1030 => x"2e8a38b4",
  1031 => x"ac5185fe",
  1032 => x"2da0fe04",
  1033 => x"bda60b80",
  1034 => x"f52d5473",
  1035 => x"80d52e09",
  1036 => x"810680ca",
  1037 => x"38bda70b",
  1038 => x"80f52d54",
  1039 => x"7381aa2e",
  1040 => x"098106ba",
  1041 => x"38800bb9",
  1042 => x"a80b80f5",
  1043 => x"2d565474",
  1044 => x"81e92e83",
  1045 => x"38815474",
  1046 => x"81eb2e8c",
  1047 => x"38805573",
  1048 => x"752e0981",
  1049 => x"0682d038",
  1050 => x"b9b30b80",
  1051 => x"f52d5574",
  1052 => x"8d38b9b4",
  1053 => x"0b80f52d",
  1054 => x"5473822e",
  1055 => x"86388055",
  1056 => x"a3b704b9",
  1057 => x"b50b80f5",
  1058 => x"2d70bfac",
  1059 => x"0cff05bf",
  1060 => x"b00cb9b6",
  1061 => x"0b80f52d",
  1062 => x"b9b70b80",
  1063 => x"f52d5876",
  1064 => x"05778280",
  1065 => x"290570bf",
  1066 => x"bc0cb9b8",
  1067 => x"0b80f52d",
  1068 => x"70bfd00c",
  1069 => x"bfb40859",
  1070 => x"57587680",
  1071 => x"2e81a338",
  1072 => x"8853b48c",
  1073 => x"52b9fa51",
  1074 => x"9cae2db8",
  1075 => x"c00881e7",
  1076 => x"38bfac08",
  1077 => x"70842bbf",
  1078 => x"b80c70bf",
  1079 => x"cc0cb9cd",
  1080 => x"0b80f52d",
  1081 => x"b9cc0b80",
  1082 => x"f52d7182",
  1083 => x"802905b9",
  1084 => x"ce0b80f5",
  1085 => x"2d708480",
  1086 => x"802912b9",
  1087 => x"cf0b80f5",
  1088 => x"2d708180",
  1089 => x"0a291270",
  1090 => x"bfd40cbf",
  1091 => x"d0087129",
  1092 => x"bfbc0805",
  1093 => x"70bfc00c",
  1094 => x"b9d50b80",
  1095 => x"f52db9d4",
  1096 => x"0b80f52d",
  1097 => x"71828029",
  1098 => x"05b9d60b",
  1099 => x"80f52d70",
  1100 => x"84808029",
  1101 => x"12b9d70b",
  1102 => x"80f52d70",
  1103 => x"982b81f0",
  1104 => x"0a067205",
  1105 => x"70bfc40c",
  1106 => x"fe117e29",
  1107 => x"7705bfc8",
  1108 => x"0c525952",
  1109 => x"43545e51",
  1110 => x"5259525d",
  1111 => x"575957a3",
  1112 => x"b004b9ba",
  1113 => x"0b80f52d",
  1114 => x"b9b90b80",
  1115 => x"f52d7182",
  1116 => x"80290570",
  1117 => x"bfb80c70",
  1118 => x"a02983ff",
  1119 => x"0570892a",
  1120 => x"70bfcc0c",
  1121 => x"b9bf0b80",
  1122 => x"f52db9be",
  1123 => x"0b80f52d",
  1124 => x"71828029",
  1125 => x"0570bfd4",
  1126 => x"0c7b7129",
  1127 => x"1e70bfc8",
  1128 => x"0c7dbfc4",
  1129 => x"0c7305bf",
  1130 => x"c00c555e",
  1131 => x"51515555",
  1132 => x"80519cec",
  1133 => x"2d815574",
  1134 => x"b8c00c02",
  1135 => x"a8050d04",
  1136 => x"02ec050d",
  1137 => x"7670872c",
  1138 => x"7180ff06",
  1139 => x"555654bf",
  1140 => x"b4088a38",
  1141 => x"73882c74",
  1142 => x"81ff0654",
  1143 => x"55b9a852",
  1144 => x"bfbc0815",
  1145 => x"519b8e2d",
  1146 => x"b8c00854",
  1147 => x"b8c00880",
  1148 => x"2eb338bf",
  1149 => x"b408802e",
  1150 => x"98387284",
  1151 => x"29b9a805",
  1152 => x"70085253",
  1153 => x"a9bc2db8",
  1154 => x"c008f00a",
  1155 => x"0653a4a3",
  1156 => x"047210b9",
  1157 => x"a8057080",
  1158 => x"e02d5253",
  1159 => x"a9ec2db8",
  1160 => x"c0085372",
  1161 => x"5473b8c0",
  1162 => x"0c029405",
  1163 => x"0d0402e0",
  1164 => x"050d7970",
  1165 => x"842cbfdc",
  1166 => x"0805718f",
  1167 => x"06525553",
  1168 => x"728938b9",
  1169 => x"a8527351",
  1170 => x"9b8e2d72",
  1171 => x"a029b9a8",
  1172 => x"05548074",
  1173 => x"80f52d56",
  1174 => x"5374732e",
  1175 => x"83388153",
  1176 => x"7481e52e",
  1177 => x"81ef3881",
  1178 => x"70740654",
  1179 => x"5872802e",
  1180 => x"81e3388b",
  1181 => x"1480f52d",
  1182 => x"70832a79",
  1183 => x"06585676",
  1184 => x"9838b784",
  1185 => x"08537288",
  1186 => x"3872bda8",
  1187 => x"0b81b72d",
  1188 => x"76b7840c",
  1189 => x"7353a6d7",
  1190 => x"04758f2e",
  1191 => x"09810681",
  1192 => x"b438749f",
  1193 => x"068d29bd",
  1194 => x"9b115153",
  1195 => x"811480f5",
  1196 => x"2d737081",
  1197 => x"055581b7",
  1198 => x"2d831480",
  1199 => x"f52d7370",
  1200 => x"81055581",
  1201 => x"b72d8514",
  1202 => x"80f52d73",
  1203 => x"70810555",
  1204 => x"81b72d87",
  1205 => x"1480f52d",
  1206 => x"73708105",
  1207 => x"5581b72d",
  1208 => x"891480f5",
  1209 => x"2d737081",
  1210 => x"055581b7",
  1211 => x"2d8e1480",
  1212 => x"f52d7370",
  1213 => x"81055581",
  1214 => x"b72d9014",
  1215 => x"80f52d73",
  1216 => x"70810555",
  1217 => x"81b72d92",
  1218 => x"1480f52d",
  1219 => x"73708105",
  1220 => x"5581b72d",
  1221 => x"941480f5",
  1222 => x"2d737081",
  1223 => x"055581b7",
  1224 => x"2d961480",
  1225 => x"f52d7370",
  1226 => x"81055581",
  1227 => x"b72d9814",
  1228 => x"80f52d73",
  1229 => x"70810555",
  1230 => x"81b72d9c",
  1231 => x"1480f52d",
  1232 => x"73708105",
  1233 => x"5581b72d",
  1234 => x"9e1480f5",
  1235 => x"2d7381b7",
  1236 => x"2d77b784",
  1237 => x"0c805372",
  1238 => x"b8c00c02",
  1239 => x"a0050d04",
  1240 => x"02cc050d",
  1241 => x"7e605e5a",
  1242 => x"800bbfd8",
  1243 => x"08bfdc08",
  1244 => x"595c5680",
  1245 => x"58bfb808",
  1246 => x"782e81ae",
  1247 => x"38778f06",
  1248 => x"a0175754",
  1249 => x"738f38b9",
  1250 => x"a8527651",
  1251 => x"8117579b",
  1252 => x"8e2db9a8",
  1253 => x"56807680",
  1254 => x"f52d5654",
  1255 => x"74742e83",
  1256 => x"38815474",
  1257 => x"81e52e80",
  1258 => x"f6388170",
  1259 => x"7506555c",
  1260 => x"73802e80",
  1261 => x"ea388b16",
  1262 => x"80f52d98",
  1263 => x"06597880",
  1264 => x"de388b53",
  1265 => x"7c527551",
  1266 => x"9cae2db8",
  1267 => x"c00880cf",
  1268 => x"389c1608",
  1269 => x"51a9bc2d",
  1270 => x"b8c00884",
  1271 => x"1b0c9a16",
  1272 => x"80e02d51",
  1273 => x"a9ec2db8",
  1274 => x"c008b8c0",
  1275 => x"08881c0c",
  1276 => x"b8c00855",
  1277 => x"55bfb408",
  1278 => x"802e9838",
  1279 => x"941680e0",
  1280 => x"2d51a9ec",
  1281 => x"2db8c008",
  1282 => x"902b83ff",
  1283 => x"f00a0670",
  1284 => x"16515473",
  1285 => x"881b0c78",
  1286 => x"7a0c7b54",
  1287 => x"a8e00481",
  1288 => x"1858bfb8",
  1289 => x"087826fe",
  1290 => x"d438bfb4",
  1291 => x"08802eae",
  1292 => x"387a51a3",
  1293 => x"c02db8c0",
  1294 => x"08b8c008",
  1295 => x"80ffffff",
  1296 => x"f806555b",
  1297 => x"7380ffff",
  1298 => x"fff82e92",
  1299 => x"38b8c008",
  1300 => x"fe05bfac",
  1301 => x"0829bfc0",
  1302 => x"080557a6",
  1303 => x"f3048054",
  1304 => x"73b8c00c",
  1305 => x"02b4050d",
  1306 => x"0402f405",
  1307 => x"0d747008",
  1308 => x"8105710c",
  1309 => x"7008bfb0",
  1310 => x"08065353",
  1311 => x"718e3888",
  1312 => x"130851a3",
  1313 => x"c02db8c0",
  1314 => x"0888140c",
  1315 => x"810bb8c0",
  1316 => x"0c028c05",
  1317 => x"0d0402f0",
  1318 => x"050d7588",
  1319 => x"1108fe05",
  1320 => x"bfac0829",
  1321 => x"bfc00811",
  1322 => x"7208bfb0",
  1323 => x"08060579",
  1324 => x"55535454",
  1325 => x"9b8e2d02",
  1326 => x"90050d04",
  1327 => x"02f4050d",
  1328 => x"7470882a",
  1329 => x"83fe8006",
  1330 => x"7072982a",
  1331 => x"0772882b",
  1332 => x"87fc8080",
  1333 => x"0673982b",
  1334 => x"81f00a06",
  1335 => x"71730707",
  1336 => x"b8c00c56",
  1337 => x"51535102",
  1338 => x"8c050d04",
  1339 => x"02f8050d",
  1340 => x"028e0580",
  1341 => x"f52d7488",
  1342 => x"2b077083",
  1343 => x"ffff06b8",
  1344 => x"c00c5102",
  1345 => x"88050d04",
  1346 => x"02f4050d",
  1347 => x"74767853",
  1348 => x"54528071",
  1349 => x"25973872",
  1350 => x"70810554",
  1351 => x"80f52d72",
  1352 => x"70810554",
  1353 => x"81b72dff",
  1354 => x"115170eb",
  1355 => x"38807281",
  1356 => x"b72d028c",
  1357 => x"050d0402",
  1358 => x"e8050d77",
  1359 => x"56807056",
  1360 => x"54737624",
  1361 => x"b138bfb8",
  1362 => x"08742eaa",
  1363 => x"387351a4",
  1364 => x"ae2db8c0",
  1365 => x"08b8c008",
  1366 => x"09810570",
  1367 => x"b8c00807",
  1368 => x"9f2a7705",
  1369 => x"81175757",
  1370 => x"53537476",
  1371 => x"248838bf",
  1372 => x"b8087426",
  1373 => x"d83872b8",
  1374 => x"c00c0298",
  1375 => x"050d0402",
  1376 => x"f0050db8",
  1377 => x"bc081651",
  1378 => x"aab72db8",
  1379 => x"c008802e",
  1380 => x"9b388b53",
  1381 => x"b8c00852",
  1382 => x"bda851aa",
  1383 => x"882dbfe4",
  1384 => x"08547380",
  1385 => x"2e8638bd",
  1386 => x"a851732d",
  1387 => x"0290050d",
  1388 => x"0402dc05",
  1389 => x"0d80705a",
  1390 => x"5574b8bc",
  1391 => x"0825af38",
  1392 => x"bfb80875",
  1393 => x"2ea83878",
  1394 => x"51a4ae2d",
  1395 => x"b8c00809",
  1396 => x"810570b8",
  1397 => x"c008079f",
  1398 => x"2a760581",
  1399 => x"1b5b5654",
  1400 => x"74b8bc08",
  1401 => x"258838bf",
  1402 => x"b8087926",
  1403 => x"da388055",
  1404 => x"78bfb808",
  1405 => x"2781cd38",
  1406 => x"7851a4ae",
  1407 => x"2db8c008",
  1408 => x"802e81a2",
  1409 => x"38b8c008",
  1410 => x"8b0580f5",
  1411 => x"2d70842a",
  1412 => x"70810677",
  1413 => x"1078842b",
  1414 => x"bda80b80",
  1415 => x"f52d5c5c",
  1416 => x"53515556",
  1417 => x"73802e80",
  1418 => x"c6387416",
  1419 => x"822bade7",
  1420 => x"0bb79012",
  1421 => x"0c547775",
  1422 => x"3110bfe8",
  1423 => x"11555690",
  1424 => x"74708105",
  1425 => x"5681b72d",
  1426 => x"a07481b7",
  1427 => x"2d7681ff",
  1428 => x"06811658",
  1429 => x"5473802e",
  1430 => x"89389c53",
  1431 => x"bda852ac",
  1432 => x"e8048b53",
  1433 => x"b8c00852",
  1434 => x"bfea1651",
  1435 => x"ad9e0474",
  1436 => x"16822baa",
  1437 => x"ff0bb790",
  1438 => x"120c5476",
  1439 => x"81ff0681",
  1440 => x"16585473",
  1441 => x"802e8938",
  1442 => x"9c53bda8",
  1443 => x"52ad9604",
  1444 => x"8b53b8c0",
  1445 => x"08527775",
  1446 => x"3110bfe8",
  1447 => x"05517655",
  1448 => x"aa882dad",
  1449 => x"b9047490",
  1450 => x"29753170",
  1451 => x"10bfe805",
  1452 => x"5154b8c0",
  1453 => x"087481b7",
  1454 => x"2d811959",
  1455 => x"748b24a2",
  1456 => x"38abf004",
  1457 => x"74902975",
  1458 => x"317010bf",
  1459 => x"e8058c77",
  1460 => x"31575154",
  1461 => x"807481b7",
  1462 => x"2d9e14ff",
  1463 => x"16565474",
  1464 => x"f33802a4",
  1465 => x"050d0402",
  1466 => x"fc050db8",
  1467 => x"bc081351",
  1468 => x"aab72db8",
  1469 => x"c008802e",
  1470 => x"8838b8c0",
  1471 => x"08519cec",
  1472 => x"2d800bb8",
  1473 => x"bc0cabb1",
  1474 => x"2d8ea32d",
  1475 => x"0284050d",
  1476 => x"0402fc05",
  1477 => x"0d725170",
  1478 => x"fd2ead38",
  1479 => x"70fd248a",
  1480 => x"3870fc2e",
  1481 => x"80c438ae",
  1482 => x"f20470fe",
  1483 => x"2eb13870",
  1484 => x"ff2e0981",
  1485 => x"06bc38b8",
  1486 => x"bc085170",
  1487 => x"802eb338",
  1488 => x"ff11b8bc",
  1489 => x"0caef204",
  1490 => x"b8bc08f0",
  1491 => x"0570b8bc",
  1492 => x"0c517080",
  1493 => x"259c3880",
  1494 => x"0bb8bc0c",
  1495 => x"aef204b8",
  1496 => x"bc088105",
  1497 => x"b8bc0cae",
  1498 => x"f204b8bc",
  1499 => x"089005b8",
  1500 => x"bc0cabb1",
  1501 => x"2d8ea32d",
  1502 => x"0284050d",
  1503 => x"0402fc05",
  1504 => x"0d800bb8",
  1505 => x"bc0cabb1",
  1506 => x"2d8dba2d",
  1507 => x"b8c008b8",
  1508 => x"ac0cb788",
  1509 => x"518fbe2d",
  1510 => x"0284050d",
  1511 => x"0471bfe4",
  1512 => x"0c040000",
  1513 => x"00ffffff",
  1514 => x"ff00ffff",
  1515 => x"ffff00ff",
  1516 => x"ffffff00",
  1517 => x"20203d56",
  1518 => x"6964656f",
  1519 => x"7061632f",
  1520 => x"4f646479",
  1521 => x"73657932",
  1522 => x"3d202000",
  1523 => x"20202020",
  1524 => x"20202020",
  1525 => x"20202020",
  1526 => x"20202020",
  1527 => x"20202020",
  1528 => x"20202000",
  1529 => x"52657365",
  1530 => x"74000000",
  1531 => x"43617267",
  1532 => x"61722043",
  1533 => x"61727475",
  1534 => x"63686f2f",
  1535 => x"466f6e74",
  1536 => x"20100000",
  1537 => x"45786974",
  1538 => x"00000000",
  1539 => x"53797374",
  1540 => x"656d3a20",
  1541 => x"4f647973",
  1542 => x"73657932",
  1543 => x"00000000",
  1544 => x"53797374",
  1545 => x"656d3a20",
  1546 => x"56696465",
  1547 => x"6f706163",
  1548 => x"00000000",
  1549 => x"47373230",
  1550 => x"30204d6f",
  1551 => x"64653a20",
  1552 => x"4f666600",
  1553 => x"47373230",
  1554 => x"30204d6f",
  1555 => x"64653a20",
  1556 => x"436f6e74",
  1557 => x"72617374",
  1558 => x"20310000",
  1559 => x"47373230",
  1560 => x"30204d6f",
  1561 => x"64653a20",
  1562 => x"436f6e74",
  1563 => x"72617374",
  1564 => x"20320000",
  1565 => x"47373230",
  1566 => x"30204d6f",
  1567 => x"64653a20",
  1568 => x"436f6e74",
  1569 => x"72617374",
  1570 => x"20330000",
  1571 => x"47373230",
  1572 => x"30204d6f",
  1573 => x"64653a20",
  1574 => x"436f6e74",
  1575 => x"72617374",
  1576 => x"20340000",
  1577 => x"47373230",
  1578 => x"30204d6f",
  1579 => x"64653a20",
  1580 => x"436f6e74",
  1581 => x"72617374",
  1582 => x"20350000",
  1583 => x"47373230",
  1584 => x"30204d6f",
  1585 => x"64653a20",
  1586 => x"436f6e74",
  1587 => x"72617374",
  1588 => x"20360000",
  1589 => x"47373230",
  1590 => x"30204d6f",
  1591 => x"64653a20",
  1592 => x"436f6e74",
  1593 => x"72617374",
  1594 => x"20370000",
  1595 => x"54686520",
  1596 => x"566f6963",
  1597 => x"653a204f",
  1598 => x"66660000",
  1599 => x"54686520",
  1600 => x"566f6963",
  1601 => x"653a204f",
  1602 => x"6e000000",
  1603 => x"53776170",
  1604 => x"204a6f79",
  1605 => x"3a204f66",
  1606 => x"66000000",
  1607 => x"53776170",
  1608 => x"206a6f79",
  1609 => x"3a204f6e",
  1610 => x"00000000",
  1611 => x"5363616e",
  1612 => x"6c696e65",
  1613 => x"733a204e",
  1614 => x"6f6e6500",
  1615 => x"5363616e",
  1616 => x"6c696e65",
  1617 => x"733a2043",
  1618 => x"52542032",
  1619 => x"35250000",
  1620 => x"5363616e",
  1621 => x"6c696e65",
  1622 => x"733a2043",
  1623 => x"52542035",
  1624 => x"30250000",
  1625 => x"5363616e",
  1626 => x"6c696e65",
  1627 => x"733a2043",
  1628 => x"52542037",
  1629 => x"35250000",
  1630 => x"43617267",
  1631 => x"61204661",
  1632 => x"6c6c6964",
  1633 => x"61000000",
  1634 => x"4f4b0000",
  1635 => x"16200000",
  1636 => x"14200000",
  1637 => x"15200000",
  1638 => x"53442069",
  1639 => x"6e69742e",
  1640 => x"2e2e0a00",
  1641 => x"53442063",
  1642 => x"61726420",
  1643 => x"72657365",
  1644 => x"74206661",
  1645 => x"696c6564",
  1646 => x"210a0000",
  1647 => x"53444843",
  1648 => x"20657272",
  1649 => x"6f72210a",
  1650 => x"00000000",
  1651 => x"57726974",
  1652 => x"65206661",
  1653 => x"696c6564",
  1654 => x"0a000000",
  1655 => x"52656164",
  1656 => x"20666169",
  1657 => x"6c65640a",
  1658 => x"00000000",
  1659 => x"43617264",
  1660 => x"20696e69",
  1661 => x"74206661",
  1662 => x"696c6564",
  1663 => x"0a000000",
  1664 => x"46415431",
  1665 => x"36202020",
  1666 => x"00000000",
  1667 => x"46415433",
  1668 => x"32202020",
  1669 => x"00000000",
  1670 => x"4e6f2070",
  1671 => x"61727469",
  1672 => x"74696f6e",
  1673 => x"20736967",
  1674 => x"0a000000",
  1675 => x"42616420",
  1676 => x"70617274",
  1677 => x"0a000000",
  1678 => x"4261636b",
  1679 => x"00000000",
  1680 => x"00000002",
  1681 => x"00000002",
  1682 => x"000017b4",
  1683 => x"00000000",
  1684 => x"00000002",
  1685 => x"000017cc",
  1686 => x"00000000",
  1687 => x"00000002",
  1688 => x"000017e4",
  1689 => x"0000034e",
  1690 => x"00000003",
  1691 => x"00001b00",
  1692 => x"00000004",
  1693 => x"00000003",
  1694 => x"00001af8",
  1695 => x"00000002",
  1696 => x"00000003",
  1697 => x"00001af0",
  1698 => x"00000002",
  1699 => x"00000003",
  1700 => x"00001ad0",
  1701 => x"00000008",
  1702 => x"00000003",
  1703 => x"00001ac8",
  1704 => x"00000002",
  1705 => x"00000002",
  1706 => x"000017ec",
  1707 => x"0000177d",
  1708 => x"00000002",
  1709 => x"00001804",
  1710 => x"000006c1",
  1711 => x"00000000",
  1712 => x"00000000",
  1713 => x"00000000",
  1714 => x"0000180c",
  1715 => x"00001820",
  1716 => x"00001834",
  1717 => x"00001844",
  1718 => x"0000185c",
  1719 => x"00001874",
  1720 => x"0000188c",
  1721 => x"000018a4",
  1722 => x"000018bc",
  1723 => x"000018d4",
  1724 => x"000018ec",
  1725 => x"000018fc",
  1726 => x"0000190c",
  1727 => x"0000191c",
  1728 => x"0000192c",
  1729 => x"0000193c",
  1730 => x"00001950",
  1731 => x"00001964",
  1732 => x"00000004",
  1733 => x"00001978",
  1734 => x"00001b10",
  1735 => x"00000004",
  1736 => x"00001988",
  1737 => x"00001a44",
  1738 => x"00000000",
  1739 => x"00000000",
  1740 => x"00000000",
  1741 => x"00000000",
  1742 => x"00000000",
  1743 => x"00000000",
  1744 => x"00000000",
  1745 => x"00000000",
  1746 => x"00000000",
  1747 => x"00000000",
  1748 => x"00000000",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"00000000",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000000",
  1755 => x"00000000",
  1756 => x"00000000",
  1757 => x"00000000",
  1758 => x"00000000",
  1759 => x"00000000",
  1760 => x"00000000",
  1761 => x"00000000",
  1762 => x"00000002",
  1763 => x"00001fe8",
  1764 => x"0000157f",
  1765 => x"00000002",
  1766 => x"00002006",
  1767 => x"0000157f",
  1768 => x"00000002",
  1769 => x"00002024",
  1770 => x"0000157f",
  1771 => x"00000002",
  1772 => x"00002042",
  1773 => x"0000157f",
  1774 => x"00000002",
  1775 => x"00002060",
  1776 => x"0000157f",
  1777 => x"00000002",
  1778 => x"0000207e",
  1779 => x"0000157f",
  1780 => x"00000002",
  1781 => x"0000209c",
  1782 => x"0000157f",
  1783 => x"00000002",
  1784 => x"000020ba",
  1785 => x"0000157f",
  1786 => x"00000002",
  1787 => x"000020d8",
  1788 => x"0000157f",
  1789 => x"00000002",
  1790 => x"000020f6",
  1791 => x"0000157f",
  1792 => x"00000002",
  1793 => x"00002114",
  1794 => x"0000157f",
  1795 => x"00000002",
  1796 => x"00002132",
  1797 => x"0000157f",
  1798 => x"00000002",
  1799 => x"00002150",
  1800 => x"0000157f",
  1801 => x"00000004",
  1802 => x"00001a38",
  1803 => x"00000000",
  1804 => x"00000000",
  1805 => x"00000000",
  1806 => x"00001711",
  1807 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

