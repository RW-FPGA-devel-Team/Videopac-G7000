-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bb6",
     9 => x"e4080b0b",
    10 => x"0bb6e808",
    11 => x"0b0b0bb6",
    12 => x"ec080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"b6ec0c0b",
    16 => x"0b0bb6e8",
    17 => x"0c0b0b0b",
    18 => x"b6e40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bafa0",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"b6e47080",
    57 => x"c194278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e604",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bb6f40c",
    65 => x"9f0bb6f8",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"b6f808ff",
    69 => x"05b6f80c",
    70 => x"b6f80880",
    71 => x"25eb38b6",
    72 => x"f408ff05",
    73 => x"b6f40cb6",
    74 => x"f4088025",
    75 => x"d738800b",
    76 => x"b6f80c80",
    77 => x"0bb6f40c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bb6f408",
    97 => x"258f3882",
    98 => x"bd2db6f4",
    99 => x"08ff05b6",
   100 => x"f40c82ff",
   101 => x"04b6f408",
   102 => x"b6f80853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"b6f408a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134b6f8",
   111 => x"088105b6",
   112 => x"f80cb6f8",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bb6f80c",
   116 => x"b6f40881",
   117 => x"05b6f40c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134b6",
   122 => x"f8088105",
   123 => x"b6f80cb6",
   124 => x"f808a02e",
   125 => x"0981068e",
   126 => x"38800bb6",
   127 => x"f80cb6f4",
   128 => x"088105b6",
   129 => x"f40c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bb6fc",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bb6fc0c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872b6",
   169 => x"fc088407",
   170 => x"b6fc0c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb2fc",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"b6fc0852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"b6e40c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c8dbf2d",
   216 => x"0284050d",
   217 => x"0402fc05",
   218 => x"0dec5192",
   219 => x"710c86a4",
   220 => x"2d82710c",
   221 => x"0284050d",
   222 => x"0402d005",
   223 => x"0d7d5480",
   224 => x"5ba40bec",
   225 => x"0c7352b7",
   226 => x"8051a6de",
   227 => x"2db6e408",
   228 => x"7b2e81ab",
   229 => x"38b78408",
   230 => x"70f80c89",
   231 => x"1580f52d",
   232 => x"8a1680f5",
   233 => x"2d718280",
   234 => x"29058817",
   235 => x"80f52d70",
   236 => x"84808029",
   237 => x"12f40c7e",
   238 => x"ff155c5e",
   239 => x"57555658",
   240 => x"767b2e8b",
   241 => x"38811a77",
   242 => x"812a585a",
   243 => x"76f738f7",
   244 => x"1a5a815b",
   245 => x"80782580",
   246 => x"e6387952",
   247 => x"7651848b",
   248 => x"2db7cc52",
   249 => x"b78051a9",
   250 => x"942db6e4",
   251 => x"08802eb8",
   252 => x"38b7cc5c",
   253 => x"83fc597b",
   254 => x"7084055d",
   255 => x"087081ff",
   256 => x"0671882a",
   257 => x"7081ff06",
   258 => x"73902a70",
   259 => x"81ff0675",
   260 => x"982ae80c",
   261 => x"e80c58e8",
   262 => x"0c57e80c",
   263 => x"fc1a5a53",
   264 => x"788025d3",
   265 => x"3888af04",
   266 => x"b6e4085b",
   267 => x"848058b7",
   268 => x"8051a8e7",
   269 => x"2dfc8018",
   270 => x"81185858",
   271 => x"87d40486",
   272 => x"b72d800b",
   273 => x"ec0c7a80",
   274 => x"2e8d38b3",
   275 => x"80518fbc",
   276 => x"2d8dbf2d",
   277 => x"88dd04b4",
   278 => x"b4518fbc",
   279 => x"2d7ab6e4",
   280 => x"0c02b005",
   281 => x"0d0402ec",
   282 => x"050d850b",
   283 => x"ec0c8da0",
   284 => x"2d8a8a2d",
   285 => x"81f82d9d",
   286 => x"fb2db6e4",
   287 => x"08802e80",
   288 => x"f43886f9",
   289 => x"51af9b2d",
   290 => x"b380518f",
   291 => x"bc2d8dbf",
   292 => x"2d8a962d",
   293 => x"8fcc2db3",
   294 => x"b80b80f5",
   295 => x"2d70892b",
   296 => x"8c8006b3",
   297 => x"c40b80f5",
   298 => x"2d70872b",
   299 => x"818006b3",
   300 => x"d00b80f5",
   301 => x"2d701082",
   302 => x"06747307",
   303 => x"07b3dc0b",
   304 => x"80f52d70",
   305 => x"852ba006",
   306 => x"b3e80b80",
   307 => x"f52d708e",
   308 => x"2b818080",
   309 => x"06747307",
   310 => x"07fc0c54",
   311 => x"54565452",
   312 => x"57575452",
   313 => x"8652b6e4",
   314 => x"088538b6",
   315 => x"e4085271",
   316 => x"ec0c8991",
   317 => x"04800bb6",
   318 => x"e40c0294",
   319 => x"050d0471",
   320 => x"980c04ff",
   321 => x"b008b6e4",
   322 => x"0c04810b",
   323 => x"ffb00c04",
   324 => x"800bffb0",
   325 => x"0c0402f4",
   326 => x"050d8b98",
   327 => x"04b6e408",
   328 => x"81f02e09",
   329 => x"81068938",
   330 => x"810bb598",
   331 => x"0c8b9804",
   332 => x"b6e40881",
   333 => x"e02e0981",
   334 => x"06893881",
   335 => x"0bb59c0c",
   336 => x"8b9804b6",
   337 => x"e40852b5",
   338 => x"9c08802e",
   339 => x"8838b6e4",
   340 => x"08818005",
   341 => x"5271842c",
   342 => x"728f0653",
   343 => x"53b59808",
   344 => x"802e9938",
   345 => x"728429b4",
   346 => x"d8057213",
   347 => x"81712b70",
   348 => x"09730806",
   349 => x"730c5153",
   350 => x"538b8e04",
   351 => x"728429b4",
   352 => x"d8057213",
   353 => x"83712b72",
   354 => x"0807720c",
   355 => x"5353800b",
   356 => x"b59c0c80",
   357 => x"0bb5980c",
   358 => x"b78c518c",
   359 => x"992db6e4",
   360 => x"08ff24fe",
   361 => x"f838800b",
   362 => x"b6e40c02",
   363 => x"8c050d04",
   364 => x"02f8050d",
   365 => x"b4d8528f",
   366 => x"51807270",
   367 => x"8405540c",
   368 => x"ff115170",
   369 => x"8025f238",
   370 => x"0288050d",
   371 => x"0402f005",
   372 => x"0d75518a",
   373 => x"902d7082",
   374 => x"2cfc06b4",
   375 => x"d8117210",
   376 => x"9e067108",
   377 => x"70722a70",
   378 => x"83068274",
   379 => x"2b700974",
   380 => x"06760c54",
   381 => x"51565753",
   382 => x"51538a8a",
   383 => x"2d71b6e4",
   384 => x"0c029005",
   385 => x"0d0402fc",
   386 => x"050d7251",
   387 => x"80710c80",
   388 => x"0b84120c",
   389 => x"0284050d",
   390 => x"0402f005",
   391 => x"0d757008",
   392 => x"84120853",
   393 => x"5353ff54",
   394 => x"71712ea8",
   395 => x"388a902d",
   396 => x"84130870",
   397 => x"84291488",
   398 => x"11700870",
   399 => x"81ff0684",
   400 => x"18088111",
   401 => x"8706841a",
   402 => x"0c535155",
   403 => x"5151518a",
   404 => x"8a2d7154",
   405 => x"73b6e40c",
   406 => x"0290050d",
   407 => x"0402f805",
   408 => x"0d8a902d",
   409 => x"e008708b",
   410 => x"2a708106",
   411 => x"51525270",
   412 => x"802e9d38",
   413 => x"b78c0870",
   414 => x"8429b794",
   415 => x"057381ff",
   416 => x"06710c51",
   417 => x"51b78c08",
   418 => x"81118706",
   419 => x"b78c0c51",
   420 => x"800bb7b4",
   421 => x"0c8a832d",
   422 => x"8a8a2d02",
   423 => x"88050d04",
   424 => x"02fc050d",
   425 => x"b78c518c",
   426 => x"862d8bb0",
   427 => x"2d8cdd51",
   428 => x"89ff2d02",
   429 => x"84050d04",
   430 => x"b7b808b6",
   431 => x"e40c0402",
   432 => x"fc050d8d",
   433 => x"c9048a96",
   434 => x"2d80f651",
   435 => x"8bcd2db6",
   436 => x"e408f338",
   437 => x"80da518b",
   438 => x"cd2db6e4",
   439 => x"08e838b6",
   440 => x"e408b5a4",
   441 => x"0cb6e408",
   442 => x"5184f02d",
   443 => x"0284050d",
   444 => x"0402ec05",
   445 => x"0d765480",
   446 => x"52870b88",
   447 => x"1580f52d",
   448 => x"56537472",
   449 => x"248338a0",
   450 => x"53725182",
   451 => x"f92d8112",
   452 => x"8b1580f5",
   453 => x"2d545272",
   454 => x"7225de38",
   455 => x"0294050d",
   456 => x"0402f005",
   457 => x"0db7b808",
   458 => x"5481f82d",
   459 => x"800bb7bc",
   460 => x"0c730880",
   461 => x"2e818038",
   462 => x"820bb6f8",
   463 => x"0cb7bc08",
   464 => x"8f06b6f4",
   465 => x"0c730852",
   466 => x"71832e96",
   467 => x"38718326",
   468 => x"89387181",
   469 => x"2eaf388f",
   470 => x"a2047185",
   471 => x"2e9f388f",
   472 => x"a2048814",
   473 => x"80f52d84",
   474 => x"1508b1c8",
   475 => x"53545285",
   476 => x"fe2d7184",
   477 => x"29137008",
   478 => x"52528fa6",
   479 => x"0473518d",
   480 => x"f12d8fa2",
   481 => x"04b5a008",
   482 => x"8815082c",
   483 => x"70810651",
   484 => x"5271802e",
   485 => x"8738b1cc",
   486 => x"518f9f04",
   487 => x"b1d05185",
   488 => x"fe2d8414",
   489 => x"085185fe",
   490 => x"2db7bc08",
   491 => x"8105b7bc",
   492 => x"0c8c1454",
   493 => x"8eb10402",
   494 => x"90050d04",
   495 => x"71b7b80c",
   496 => x"8ea12db7",
   497 => x"bc08ff05",
   498 => x"b7c00c04",
   499 => x"02e8050d",
   500 => x"b7b808b7",
   501 => x"c4085755",
   502 => x"87518bcd",
   503 => x"2db6e408",
   504 => x"812a7081",
   505 => x"06515271",
   506 => x"802ea038",
   507 => x"8ff2048a",
   508 => x"962d8751",
   509 => x"8bcd2db6",
   510 => x"e408f438",
   511 => x"b5a40881",
   512 => x"3270b5a4",
   513 => x"0c705252",
   514 => x"84f02d80",
   515 => x"fe518bcd",
   516 => x"2db6e408",
   517 => x"802ea638",
   518 => x"b5a40880",
   519 => x"2e913880",
   520 => x"0bb5a40c",
   521 => x"805184f0",
   522 => x"2d90af04",
   523 => x"8a962d80",
   524 => x"fe518bcd",
   525 => x"2db6e408",
   526 => x"f33886e5",
   527 => x"2db5a408",
   528 => x"903881fd",
   529 => x"518bcd2d",
   530 => x"81fa518b",
   531 => x"cd2d9682",
   532 => x"0481f551",
   533 => x"8bcd2db6",
   534 => x"e408812a",
   535 => x"70810651",
   536 => x"5271802e",
   537 => x"af38b7c0",
   538 => x"08527180",
   539 => x"2e8938ff",
   540 => x"12b7c00c",
   541 => x"919404b7",
   542 => x"bc0810b7",
   543 => x"bc080570",
   544 => x"84291651",
   545 => x"52881208",
   546 => x"802e8938",
   547 => x"ff518812",
   548 => x"0852712d",
   549 => x"81f2518b",
   550 => x"cd2db6e4",
   551 => x"08812a70",
   552 => x"81065152",
   553 => x"71802eb1",
   554 => x"38b7bc08",
   555 => x"ff11b7c0",
   556 => x"08565353",
   557 => x"73722589",
   558 => x"388114b7",
   559 => x"c00c91d9",
   560 => x"04721013",
   561 => x"70842916",
   562 => x"51528812",
   563 => x"08802e89",
   564 => x"38fe5188",
   565 => x"12085271",
   566 => x"2d81fd51",
   567 => x"8bcd2db6",
   568 => x"e408812a",
   569 => x"70810651",
   570 => x"5271802e",
   571 => x"ad38b7c0",
   572 => x"08802e89",
   573 => x"38800bb7",
   574 => x"c00c929a",
   575 => x"04b7bc08",
   576 => x"10b7bc08",
   577 => x"05708429",
   578 => x"16515288",
   579 => x"1208802e",
   580 => x"8938fd51",
   581 => x"88120852",
   582 => x"712d81fa",
   583 => x"518bcd2d",
   584 => x"b6e40881",
   585 => x"2a708106",
   586 => x"51527180",
   587 => x"2eae38b7",
   588 => x"bc08ff11",
   589 => x"5452b7c0",
   590 => x"08732588",
   591 => x"3872b7c0",
   592 => x"0c92dc04",
   593 => x"71101270",
   594 => x"84291651",
   595 => x"52881208",
   596 => x"802e8938",
   597 => x"fc518812",
   598 => x"0852712d",
   599 => x"b7c00870",
   600 => x"53547380",
   601 => x"2e8a388c",
   602 => x"15ff1555",
   603 => x"5592e204",
   604 => x"820bb6f8",
   605 => x"0c718f06",
   606 => x"b6f40c81",
   607 => x"eb518bcd",
   608 => x"2db6e408",
   609 => x"812a7081",
   610 => x"06515271",
   611 => x"802ead38",
   612 => x"7408852e",
   613 => x"098106a4",
   614 => x"38881580",
   615 => x"f52dff05",
   616 => x"52718816",
   617 => x"81b72d71",
   618 => x"982b5271",
   619 => x"80258838",
   620 => x"800b8816",
   621 => x"81b72d74",
   622 => x"518df12d",
   623 => x"81f4518b",
   624 => x"cd2db6e4",
   625 => x"08812a70",
   626 => x"81065152",
   627 => x"71802eb3",
   628 => x"38740885",
   629 => x"2e098106",
   630 => x"aa388815",
   631 => x"80f52d81",
   632 => x"05527188",
   633 => x"1681b72d",
   634 => x"7181ff06",
   635 => x"8b1680f5",
   636 => x"2d545272",
   637 => x"72278738",
   638 => x"72881681",
   639 => x"b72d7451",
   640 => x"8df12d80",
   641 => x"da518bcd",
   642 => x"2db6e408",
   643 => x"812a7081",
   644 => x"06515271",
   645 => x"802e81a6",
   646 => x"38b7b808",
   647 => x"b7c00855",
   648 => x"5373802e",
   649 => x"8a388c13",
   650 => x"ff155553",
   651 => x"94a10472",
   652 => x"08527182",
   653 => x"2ea63871",
   654 => x"82268938",
   655 => x"71812ea9",
   656 => x"3895be04",
   657 => x"71832eb1",
   658 => x"3871842e",
   659 => x"09810680",
   660 => x"ed388813",
   661 => x"08518fbc",
   662 => x"2d95be04",
   663 => x"b7c00851",
   664 => x"88130852",
   665 => x"712d95be",
   666 => x"04810b88",
   667 => x"14082bb5",
   668 => x"a00832b5",
   669 => x"a00c9594",
   670 => x"04881380",
   671 => x"f52d8105",
   672 => x"8b1480f5",
   673 => x"2d535471",
   674 => x"74248338",
   675 => x"80547388",
   676 => x"1481b72d",
   677 => x"8ea12d95",
   678 => x"be047508",
   679 => x"802ea238",
   680 => x"7508518b",
   681 => x"cd2db6e4",
   682 => x"08810652",
   683 => x"71802e8b",
   684 => x"38b7c008",
   685 => x"51841608",
   686 => x"52712d88",
   687 => x"165675da",
   688 => x"38805480",
   689 => x"0bb6f80c",
   690 => x"738f06b6",
   691 => x"f40ca052",
   692 => x"73b7c008",
   693 => x"2e098106",
   694 => x"9838b7bc",
   695 => x"08ff0574",
   696 => x"32700981",
   697 => x"05707207",
   698 => x"9f2a9171",
   699 => x"31515153",
   700 => x"53715182",
   701 => x"f92d8114",
   702 => x"548e7425",
   703 => x"c638b5a4",
   704 => x"085271b6",
   705 => x"e40c0298",
   706 => x"050d0402",
   707 => x"f4050dd4",
   708 => x"5281ff72",
   709 => x"0c710853",
   710 => x"81ff720c",
   711 => x"72882b83",
   712 => x"fe800672",
   713 => x"087081ff",
   714 => x"06515253",
   715 => x"81ff720c",
   716 => x"72710788",
   717 => x"2b720870",
   718 => x"81ff0651",
   719 => x"525381ff",
   720 => x"720c7271",
   721 => x"07882b72",
   722 => x"087081ff",
   723 => x"067207b6",
   724 => x"e40c5253",
   725 => x"028c050d",
   726 => x"0402f405",
   727 => x"0d747671",
   728 => x"81ff06d4",
   729 => x"0c5353b7",
   730 => x"c8088538",
   731 => x"71892b52",
   732 => x"71982ad4",
   733 => x"0c71902a",
   734 => x"7081ff06",
   735 => x"d40c5171",
   736 => x"882a7081",
   737 => x"ff06d40c",
   738 => x"517181ff",
   739 => x"06d40c72",
   740 => x"902a7081",
   741 => x"ff06d40c",
   742 => x"51d40870",
   743 => x"81ff0651",
   744 => x"5182b8bf",
   745 => x"527081ff",
   746 => x"2e098106",
   747 => x"943881ff",
   748 => x"0bd40cd4",
   749 => x"087081ff",
   750 => x"06ff1454",
   751 => x"515171e5",
   752 => x"3870b6e4",
   753 => x"0c028c05",
   754 => x"0d0402fc",
   755 => x"050d81c7",
   756 => x"5181ff0b",
   757 => x"d40cff11",
   758 => x"51708025",
   759 => x"f4380284",
   760 => x"050d0402",
   761 => x"f4050d81",
   762 => x"ff0bd40c",
   763 => x"93538052",
   764 => x"87fc80c1",
   765 => x"5196d92d",
   766 => x"b6e4088b",
   767 => x"3881ff0b",
   768 => x"d40c8153",
   769 => x"98900497",
   770 => x"ca2dff13",
   771 => x"5372df38",
   772 => x"72b6e40c",
   773 => x"028c050d",
   774 => x"0402ec05",
   775 => x"0d810bb7",
   776 => x"c80c8454",
   777 => x"d008708f",
   778 => x"2a708106",
   779 => x"51515372",
   780 => x"f33872d0",
   781 => x"0c97ca2d",
   782 => x"b1d45185",
   783 => x"fe2dd008",
   784 => x"708f2a70",
   785 => x"81065151",
   786 => x"5372f338",
   787 => x"810bd00c",
   788 => x"b1538052",
   789 => x"84d480c0",
   790 => x"5196d92d",
   791 => x"b6e40881",
   792 => x"2e933872",
   793 => x"822ebd38",
   794 => x"ff135372",
   795 => x"e538ff14",
   796 => x"5473ffb0",
   797 => x"3897ca2d",
   798 => x"83aa5284",
   799 => x"9c80c851",
   800 => x"96d92db6",
   801 => x"e408812e",
   802 => x"09810692",
   803 => x"38968b2d",
   804 => x"b6e40883",
   805 => x"ffff0653",
   806 => x"7283aa2e",
   807 => x"9d3897e3",
   808 => x"2d99b504",
   809 => x"b1e05185",
   810 => x"fe2d8053",
   811 => x"9b8304b1",
   812 => x"f85185fe",
   813 => x"2d80549a",
   814 => x"d50481ff",
   815 => x"0bd40cb1",
   816 => x"5497ca2d",
   817 => x"8fcf5380",
   818 => x"5287fc80",
   819 => x"f75196d9",
   820 => x"2db6e408",
   821 => x"55b6e408",
   822 => x"812e0981",
   823 => x"069b3881",
   824 => x"ff0bd40c",
   825 => x"820a5284",
   826 => x"9c80e951",
   827 => x"96d92db6",
   828 => x"e408802e",
   829 => x"8d3897ca",
   830 => x"2dff1353",
   831 => x"72c9389a",
   832 => x"c80481ff",
   833 => x"0bd40cb6",
   834 => x"e4085287",
   835 => x"fc80fa51",
   836 => x"96d92db6",
   837 => x"e408b138",
   838 => x"81ff0bd4",
   839 => x"0cd40853",
   840 => x"81ff0bd4",
   841 => x"0c81ff0b",
   842 => x"d40c81ff",
   843 => x"0bd40c81",
   844 => x"ff0bd40c",
   845 => x"72862a70",
   846 => x"81067656",
   847 => x"51537295",
   848 => x"38b6e408",
   849 => x"549ad504",
   850 => x"73822efe",
   851 => x"e238ff14",
   852 => x"5473feed",
   853 => x"3873b7c8",
   854 => x"0c738b38",
   855 => x"815287fc",
   856 => x"80d05196",
   857 => x"d92d81ff",
   858 => x"0bd40cd0",
   859 => x"08708f2a",
   860 => x"70810651",
   861 => x"515372f3",
   862 => x"3872d00c",
   863 => x"81ff0bd4",
   864 => x"0c815372",
   865 => x"b6e40c02",
   866 => x"94050d04",
   867 => x"02e8050d",
   868 => x"78558056",
   869 => x"81ff0bd4",
   870 => x"0cd00870",
   871 => x"8f2a7081",
   872 => x"06515153",
   873 => x"72f33882",
   874 => x"810bd00c",
   875 => x"81ff0bd4",
   876 => x"0c775287",
   877 => x"fc80d151",
   878 => x"96d92d80",
   879 => x"dbc6df54",
   880 => x"b6e40880",
   881 => x"2e8a38b2",
   882 => x"985185fe",
   883 => x"2d9ca304",
   884 => x"81ff0bd4",
   885 => x"0cd40870",
   886 => x"81ff0651",
   887 => x"537281fe",
   888 => x"2e098106",
   889 => x"9d3880ff",
   890 => x"53968b2d",
   891 => x"b6e40875",
   892 => x"70840557",
   893 => x"0cff1353",
   894 => x"728025ed",
   895 => x"3881569c",
   896 => x"8804ff14",
   897 => x"5473c938",
   898 => x"81ff0bd4",
   899 => x"0c81ff0b",
   900 => x"d40cd008",
   901 => x"708f2a70",
   902 => x"81065151",
   903 => x"5372f338",
   904 => x"72d00c75",
   905 => x"b6e40c02",
   906 => x"98050d04",
   907 => x"02e8050d",
   908 => x"77797b58",
   909 => x"55558053",
   910 => x"727625a3",
   911 => x"38747081",
   912 => x"055680f5",
   913 => x"2d747081",
   914 => x"055680f5",
   915 => x"2d525271",
   916 => x"712e8638",
   917 => x"81519ce1",
   918 => x"04811353",
   919 => x"9cb80480",
   920 => x"5170b6e4",
   921 => x"0c029805",
   922 => x"0d0402ec",
   923 => x"050d7655",
   924 => x"74802ebb",
   925 => x"389a1580",
   926 => x"e02d51a9",
   927 => x"ea2db6e4",
   928 => x"08b6e408",
   929 => x"bdfc0cb6",
   930 => x"e4085454",
   931 => x"bdd80880",
   932 => x"2e993894",
   933 => x"1580e02d",
   934 => x"51a9ea2d",
   935 => x"b6e40890",
   936 => x"2b83fff0",
   937 => x"0a067075",
   938 => x"07515372",
   939 => x"bdfc0cbd",
   940 => x"fc085372",
   941 => x"802e9938",
   942 => x"bdd008fe",
   943 => x"147129bd",
   944 => x"e40805be",
   945 => x"800c7084",
   946 => x"2bbddc0c",
   947 => x"549df604",
   948 => x"bde808bd",
   949 => x"fc0cbdec",
   950 => x"08be800c",
   951 => x"bdd80880",
   952 => x"2e8a38bd",
   953 => x"d008842b",
   954 => x"539df204",
   955 => x"bdf00884",
   956 => x"2b5372bd",
   957 => x"dc0c0294",
   958 => x"050d0402",
   959 => x"d8050d80",
   960 => x"0bbdd80c",
   961 => x"84549899",
   962 => x"2db6e408",
   963 => x"802e9538",
   964 => x"b7cc5280",
   965 => x"519b8c2d",
   966 => x"b6e40880",
   967 => x"2e8638fe",
   968 => x"549eac04",
   969 => x"ff145473",
   970 => x"8024db38",
   971 => x"738c38b2",
   972 => x"a85185fe",
   973 => x"2d7355a3",
   974 => x"b5048056",
   975 => x"810bbe84",
   976 => x"0c8853b2",
   977 => x"bc52b882",
   978 => x"519cac2d",
   979 => x"b6e40876",
   980 => x"2e098106",
   981 => x"8738b6e4",
   982 => x"08be840c",
   983 => x"8853b2c8",
   984 => x"52b89e51",
   985 => x"9cac2db6",
   986 => x"e4088738",
   987 => x"b6e408be",
   988 => x"840cbe84",
   989 => x"08802e80",
   990 => x"f638bb92",
   991 => x"0b80f52d",
   992 => x"bb930b80",
   993 => x"f52d7198",
   994 => x"2b71902b",
   995 => x"07bb940b",
   996 => x"80f52d70",
   997 => x"882b7207",
   998 => x"bb950b80",
   999 => x"f52d7107",
  1000 => x"bbca0b80",
  1001 => x"f52dbbcb",
  1002 => x"0b80f52d",
  1003 => x"71882b07",
  1004 => x"535f5452",
  1005 => x"5a565755",
  1006 => x"7381abaa",
  1007 => x"2e098106",
  1008 => x"8d387551",
  1009 => x"a9ba2db6",
  1010 => x"e408569f",
  1011 => x"db047382",
  1012 => x"d4d52e87",
  1013 => x"38b2d451",
  1014 => x"a09c04b7",
  1015 => x"cc527551",
  1016 => x"9b8c2db6",
  1017 => x"e40855b6",
  1018 => x"e408802e",
  1019 => x"83c73888",
  1020 => x"53b2c852",
  1021 => x"b89e519c",
  1022 => x"ac2db6e4",
  1023 => x"08893881",
  1024 => x"0bbdd80c",
  1025 => x"a0a20488",
  1026 => x"53b2bc52",
  1027 => x"b882519c",
  1028 => x"ac2db6e4",
  1029 => x"08802e8a",
  1030 => x"38b2e851",
  1031 => x"85fe2da0",
  1032 => x"fc04bbca",
  1033 => x"0b80f52d",
  1034 => x"547380d5",
  1035 => x"2e098106",
  1036 => x"80ca38bb",
  1037 => x"cb0b80f5",
  1038 => x"2d547381",
  1039 => x"aa2e0981",
  1040 => x"06ba3880",
  1041 => x"0bb7cc0b",
  1042 => x"80f52d56",
  1043 => x"547481e9",
  1044 => x"2e833881",
  1045 => x"547481eb",
  1046 => x"2e8c3880",
  1047 => x"5573752e",
  1048 => x"09810682",
  1049 => x"d038b7d7",
  1050 => x"0b80f52d",
  1051 => x"55748d38",
  1052 => x"b7d80b80",
  1053 => x"f52d5473",
  1054 => x"822e8638",
  1055 => x"8055a3b5",
  1056 => x"04b7d90b",
  1057 => x"80f52d70",
  1058 => x"bdd00cff",
  1059 => x"05bdd40c",
  1060 => x"b7da0b80",
  1061 => x"f52db7db",
  1062 => x"0b80f52d",
  1063 => x"58760577",
  1064 => x"82802905",
  1065 => x"70bde00c",
  1066 => x"b7dc0b80",
  1067 => x"f52d70bd",
  1068 => x"f40cbdd8",
  1069 => x"08595758",
  1070 => x"76802e81",
  1071 => x"a3388853",
  1072 => x"b2c852b8",
  1073 => x"9e519cac",
  1074 => x"2db6e408",
  1075 => x"81e738bd",
  1076 => x"d0087084",
  1077 => x"2bbddc0c",
  1078 => x"70bdf00c",
  1079 => x"b7f10b80",
  1080 => x"f52db7f0",
  1081 => x"0b80f52d",
  1082 => x"71828029",
  1083 => x"05b7f20b",
  1084 => x"80f52d70",
  1085 => x"84808029",
  1086 => x"12b7f30b",
  1087 => x"80f52d70",
  1088 => x"81800a29",
  1089 => x"1270bdf8",
  1090 => x"0cbdf408",
  1091 => x"7129bde0",
  1092 => x"080570bd",
  1093 => x"e40cb7f9",
  1094 => x"0b80f52d",
  1095 => x"b7f80b80",
  1096 => x"f52d7182",
  1097 => x"802905b7",
  1098 => x"fa0b80f5",
  1099 => x"2d708480",
  1100 => x"802912b7",
  1101 => x"fb0b80f5",
  1102 => x"2d70982b",
  1103 => x"81f00a06",
  1104 => x"720570bd",
  1105 => x"e80cfe11",
  1106 => x"7e297705",
  1107 => x"bdec0c52",
  1108 => x"59524354",
  1109 => x"5e515259",
  1110 => x"525d5759",
  1111 => x"57a3ae04",
  1112 => x"b7de0b80",
  1113 => x"f52db7dd",
  1114 => x"0b80f52d",
  1115 => x"71828029",
  1116 => x"0570bddc",
  1117 => x"0c70a029",
  1118 => x"83ff0570",
  1119 => x"892a70bd",
  1120 => x"f00cb7e3",
  1121 => x"0b80f52d",
  1122 => x"b7e20b80",
  1123 => x"f52d7182",
  1124 => x"80290570",
  1125 => x"bdf80c7b",
  1126 => x"71291e70",
  1127 => x"bdec0c7d",
  1128 => x"bde80c73",
  1129 => x"05bde40c",
  1130 => x"555e5151",
  1131 => x"55558051",
  1132 => x"9cea2d81",
  1133 => x"5574b6e4",
  1134 => x"0c02a805",
  1135 => x"0d0402ec",
  1136 => x"050d7670",
  1137 => x"872c7180",
  1138 => x"ff065556",
  1139 => x"54bdd808",
  1140 => x"8a387388",
  1141 => x"2c7481ff",
  1142 => x"065455b7",
  1143 => x"cc52bde0",
  1144 => x"0815519b",
  1145 => x"8c2db6e4",
  1146 => x"0854b6e4",
  1147 => x"08802eb3",
  1148 => x"38bdd808",
  1149 => x"802e9838",
  1150 => x"728429b7",
  1151 => x"cc057008",
  1152 => x"5253a9ba",
  1153 => x"2db6e408",
  1154 => x"f00a0653",
  1155 => x"a4a10472",
  1156 => x"10b7cc05",
  1157 => x"7080e02d",
  1158 => x"5253a9ea",
  1159 => x"2db6e408",
  1160 => x"53725473",
  1161 => x"b6e40c02",
  1162 => x"94050d04",
  1163 => x"02e0050d",
  1164 => x"7970842c",
  1165 => x"be800805",
  1166 => x"718f0652",
  1167 => x"55537289",
  1168 => x"38b7cc52",
  1169 => x"73519b8c",
  1170 => x"2d72a029",
  1171 => x"b7cc0554",
  1172 => x"807480f5",
  1173 => x"2d565374",
  1174 => x"732e8338",
  1175 => x"81537481",
  1176 => x"e52e81ef",
  1177 => x"38817074",
  1178 => x"06545872",
  1179 => x"802e81e3",
  1180 => x"388b1480",
  1181 => x"f52d7083",
  1182 => x"2a790658",
  1183 => x"56769838",
  1184 => x"b5a80853",
  1185 => x"72883872",
  1186 => x"bbcc0b81",
  1187 => x"b72d76b5",
  1188 => x"a80c7353",
  1189 => x"a6d50475",
  1190 => x"8f2e0981",
  1191 => x"0681b438",
  1192 => x"749f068d",
  1193 => x"29bbbf11",
  1194 => x"51538114",
  1195 => x"80f52d73",
  1196 => x"70810555",
  1197 => x"81b72d83",
  1198 => x"1480f52d",
  1199 => x"73708105",
  1200 => x"5581b72d",
  1201 => x"851480f5",
  1202 => x"2d737081",
  1203 => x"055581b7",
  1204 => x"2d871480",
  1205 => x"f52d7370",
  1206 => x"81055581",
  1207 => x"b72d8914",
  1208 => x"80f52d73",
  1209 => x"70810555",
  1210 => x"81b72d8e",
  1211 => x"1480f52d",
  1212 => x"73708105",
  1213 => x"5581b72d",
  1214 => x"901480f5",
  1215 => x"2d737081",
  1216 => x"055581b7",
  1217 => x"2d921480",
  1218 => x"f52d7370",
  1219 => x"81055581",
  1220 => x"b72d9414",
  1221 => x"80f52d73",
  1222 => x"70810555",
  1223 => x"81b72d96",
  1224 => x"1480f52d",
  1225 => x"73708105",
  1226 => x"5581b72d",
  1227 => x"981480f5",
  1228 => x"2d737081",
  1229 => x"055581b7",
  1230 => x"2d9c1480",
  1231 => x"f52d7370",
  1232 => x"81055581",
  1233 => x"b72d9e14",
  1234 => x"80f52d73",
  1235 => x"81b72d77",
  1236 => x"b5a80c80",
  1237 => x"5372b6e4",
  1238 => x"0c02a005",
  1239 => x"0d0402cc",
  1240 => x"050d7e60",
  1241 => x"5e5a800b",
  1242 => x"bdfc08be",
  1243 => x"8008595c",
  1244 => x"568058bd",
  1245 => x"dc08782e",
  1246 => x"81ae3877",
  1247 => x"8f06a017",
  1248 => x"5754738f",
  1249 => x"38b7cc52",
  1250 => x"76518117",
  1251 => x"579b8c2d",
  1252 => x"b7cc5680",
  1253 => x"7680f52d",
  1254 => x"56547474",
  1255 => x"2e833881",
  1256 => x"547481e5",
  1257 => x"2e80f638",
  1258 => x"81707506",
  1259 => x"555c7380",
  1260 => x"2e80ea38",
  1261 => x"8b1680f5",
  1262 => x"2d980659",
  1263 => x"7880de38",
  1264 => x"8b537c52",
  1265 => x"75519cac",
  1266 => x"2db6e408",
  1267 => x"80cf389c",
  1268 => x"160851a9",
  1269 => x"ba2db6e4",
  1270 => x"08841b0c",
  1271 => x"9a1680e0",
  1272 => x"2d51a9ea",
  1273 => x"2db6e408",
  1274 => x"b6e40888",
  1275 => x"1c0cb6e4",
  1276 => x"085555bd",
  1277 => x"d808802e",
  1278 => x"98389416",
  1279 => x"80e02d51",
  1280 => x"a9ea2db6",
  1281 => x"e408902b",
  1282 => x"83fff00a",
  1283 => x"06701651",
  1284 => x"5473881b",
  1285 => x"0c787a0c",
  1286 => x"7b54a8de",
  1287 => x"04811858",
  1288 => x"bddc0878",
  1289 => x"26fed438",
  1290 => x"bdd80880",
  1291 => x"2eae387a",
  1292 => x"51a3be2d",
  1293 => x"b6e408b6",
  1294 => x"e40880ff",
  1295 => x"fffff806",
  1296 => x"555b7380",
  1297 => x"fffffff8",
  1298 => x"2e9238b6",
  1299 => x"e408fe05",
  1300 => x"bdd00829",
  1301 => x"bde40805",
  1302 => x"57a6f104",
  1303 => x"805473b6",
  1304 => x"e40c02b4",
  1305 => x"050d0402",
  1306 => x"f4050d74",
  1307 => x"70088105",
  1308 => x"710c7008",
  1309 => x"bdd40806",
  1310 => x"5353718e",
  1311 => x"38881308",
  1312 => x"51a3be2d",
  1313 => x"b6e40888",
  1314 => x"140c810b",
  1315 => x"b6e40c02",
  1316 => x"8c050d04",
  1317 => x"02f0050d",
  1318 => x"75881108",
  1319 => x"fe05bdd0",
  1320 => x"0829bde4",
  1321 => x"08117208",
  1322 => x"bdd40806",
  1323 => x"05795553",
  1324 => x"54549b8c",
  1325 => x"2d029005",
  1326 => x"0d0402f4",
  1327 => x"050d7470",
  1328 => x"882a83fe",
  1329 => x"80067072",
  1330 => x"982a0772",
  1331 => x"882b87fc",
  1332 => x"80800673",
  1333 => x"982b81f0",
  1334 => x"0a067173",
  1335 => x"0707b6e4",
  1336 => x"0c565153",
  1337 => x"51028c05",
  1338 => x"0d0402f8",
  1339 => x"050d028e",
  1340 => x"0580f52d",
  1341 => x"74882b07",
  1342 => x"7083ffff",
  1343 => x"06b6e40c",
  1344 => x"51028805",
  1345 => x"0d0402f4",
  1346 => x"050d7476",
  1347 => x"78535452",
  1348 => x"80712597",
  1349 => x"38727081",
  1350 => x"055480f5",
  1351 => x"2d727081",
  1352 => x"055481b7",
  1353 => x"2dff1151",
  1354 => x"70eb3880",
  1355 => x"7281b72d",
  1356 => x"028c050d",
  1357 => x"0402e805",
  1358 => x"0d775680",
  1359 => x"70565473",
  1360 => x"7624b138",
  1361 => x"bddc0874",
  1362 => x"2eaa3873",
  1363 => x"51a4ac2d",
  1364 => x"b6e408b6",
  1365 => x"e4080981",
  1366 => x"0570b6e4",
  1367 => x"08079f2a",
  1368 => x"77058117",
  1369 => x"57575353",
  1370 => x"74762488",
  1371 => x"38bddc08",
  1372 => x"7426d838",
  1373 => x"72b6e40c",
  1374 => x"0298050d",
  1375 => x"0402f005",
  1376 => x"0db6e008",
  1377 => x"1651aab5",
  1378 => x"2db6e408",
  1379 => x"802e9b38",
  1380 => x"8b53b6e4",
  1381 => x"0852bbcc",
  1382 => x"51aa862d",
  1383 => x"be880854",
  1384 => x"73802e86",
  1385 => x"38bbcc51",
  1386 => x"732d0290",
  1387 => x"050d0402",
  1388 => x"dc050d80",
  1389 => x"705a5574",
  1390 => x"b6e00825",
  1391 => x"af38bddc",
  1392 => x"08752ea8",
  1393 => x"387851a4",
  1394 => x"ac2db6e4",
  1395 => x"08098105",
  1396 => x"70b6e408",
  1397 => x"079f2a76",
  1398 => x"05811b5b",
  1399 => x"565474b6",
  1400 => x"e0082588",
  1401 => x"38bddc08",
  1402 => x"7926da38",
  1403 => x"805578bd",
  1404 => x"dc082781",
  1405 => x"cd387851",
  1406 => x"a4ac2db6",
  1407 => x"e408802e",
  1408 => x"81a238b6",
  1409 => x"e4088b05",
  1410 => x"80f52d70",
  1411 => x"842a7081",
  1412 => x"06771078",
  1413 => x"842bbbcc",
  1414 => x"0b80f52d",
  1415 => x"5c5c5351",
  1416 => x"55567380",
  1417 => x"2e80c638",
  1418 => x"7416822b",
  1419 => x"ade50bb5",
  1420 => x"b4120c54",
  1421 => x"77753110",
  1422 => x"be8c1155",
  1423 => x"56907470",
  1424 => x"81055681",
  1425 => x"b72da074",
  1426 => x"81b72d76",
  1427 => x"81ff0681",
  1428 => x"16585473",
  1429 => x"802e8938",
  1430 => x"9c53bbcc",
  1431 => x"52ace604",
  1432 => x"8b53b6e4",
  1433 => x"0852be8e",
  1434 => x"1651ad9c",
  1435 => x"04741682",
  1436 => x"2baafd0b",
  1437 => x"b5b4120c",
  1438 => x"547681ff",
  1439 => x"06811658",
  1440 => x"5473802e",
  1441 => x"89389c53",
  1442 => x"bbcc52ad",
  1443 => x"94048b53",
  1444 => x"b6e40852",
  1445 => x"77753110",
  1446 => x"be8c0551",
  1447 => x"7655aa86",
  1448 => x"2dadb704",
  1449 => x"74902975",
  1450 => x"317010be",
  1451 => x"8c055154",
  1452 => x"b6e40874",
  1453 => x"81b72d81",
  1454 => x"1959748b",
  1455 => x"24a238ab",
  1456 => x"ee047490",
  1457 => x"29753170",
  1458 => x"10be8c05",
  1459 => x"8c773157",
  1460 => x"51548074",
  1461 => x"81b72d9e",
  1462 => x"14ff1656",
  1463 => x"5474f338",
  1464 => x"02a4050d",
  1465 => x"0402fc05",
  1466 => x"0db6e008",
  1467 => x"1351aab5",
  1468 => x"2db6e408",
  1469 => x"802e8838",
  1470 => x"b6e40851",
  1471 => x"9cea2d80",
  1472 => x"0bb6e00c",
  1473 => x"abaf2d8e",
  1474 => x"a12d0284",
  1475 => x"050d0402",
  1476 => x"fc050d72",
  1477 => x"5170fd2e",
  1478 => x"ad3870fd",
  1479 => x"248a3870",
  1480 => x"fc2e80c4",
  1481 => x"38aef004",
  1482 => x"70fe2eb1",
  1483 => x"3870ff2e",
  1484 => x"098106bc",
  1485 => x"38b6e008",
  1486 => x"5170802e",
  1487 => x"b338ff11",
  1488 => x"b6e00cae",
  1489 => x"f004b6e0",
  1490 => x"08f00570",
  1491 => x"b6e00c51",
  1492 => x"7080259c",
  1493 => x"38800bb6",
  1494 => x"e00caef0",
  1495 => x"04b6e008",
  1496 => x"8105b6e0",
  1497 => x"0caef004",
  1498 => x"b6e00890",
  1499 => x"05b6e00c",
  1500 => x"abaf2d8e",
  1501 => x"a12d0284",
  1502 => x"050d0402",
  1503 => x"fc050d80",
  1504 => x"0bb6e00c",
  1505 => x"abaf2d8d",
  1506 => x"b82db6e4",
  1507 => x"08b6d00c",
  1508 => x"b5ac518f",
  1509 => x"bc2d0284",
  1510 => x"050d0471",
  1511 => x"be880c04",
  1512 => x"00ffffff",
  1513 => x"ff00ffff",
  1514 => x"ffff00ff",
  1515 => x"ffffff00",
  1516 => x"2020203d",
  1517 => x"52616d70",
  1518 => x"61205669",
  1519 => x"64656f70",
  1520 => x"61633d20",
  1521 => x"20202000",
  1522 => x"20202020",
  1523 => x"20202020",
  1524 => x"20202020",
  1525 => x"20202020",
  1526 => x"20202020",
  1527 => x"20202000",
  1528 => x"52657365",
  1529 => x"74000000",
  1530 => x"43617267",
  1531 => x"61722043",
  1532 => x"61727475",
  1533 => x"63686f2f",
  1534 => x"466f6e74",
  1535 => x"20100000",
  1536 => x"45786974",
  1537 => x"00000000",
  1538 => x"4f647973",
  1539 => x"73657932",
  1540 => x"00000000",
  1541 => x"56696465",
  1542 => x"6f706163",
  1543 => x"00000000",
  1544 => x"4e747363",
  1545 => x"00000000",
  1546 => x"50616c00",
  1547 => x"54686520",
  1548 => x"566f6963",
  1549 => x"65204f66",
  1550 => x"66000000",
  1551 => x"54686520",
  1552 => x"566f6963",
  1553 => x"65204f6e",
  1554 => x"00000000",
  1555 => x"53776170",
  1556 => x"204a6f79",
  1557 => x"204f6666",
  1558 => x"00000000",
  1559 => x"53776170",
  1560 => x"206a6f79",
  1561 => x"204f6e00",
  1562 => x"5363616e",
  1563 => x"6c696e65",
  1564 => x"73204e6f",
  1565 => x"6e650000",
  1566 => x"5363616e",
  1567 => x"6c696e65",
  1568 => x"73204352",
  1569 => x"54203235",
  1570 => x"25000000",
  1571 => x"5363616e",
  1572 => x"6c696e65",
  1573 => x"73204352",
  1574 => x"54203530",
  1575 => x"25000000",
  1576 => x"5363616e",
  1577 => x"6c696e65",
  1578 => x"73204352",
  1579 => x"54203735",
  1580 => x"25000000",
  1581 => x"43617267",
  1582 => x"61204661",
  1583 => x"6c6c6964",
  1584 => x"61000000",
  1585 => x"4f4b0000",
  1586 => x"16200000",
  1587 => x"14200000",
  1588 => x"15200000",
  1589 => x"53442069",
  1590 => x"6e69742e",
  1591 => x"2e2e0a00",
  1592 => x"53442063",
  1593 => x"61726420",
  1594 => x"72657365",
  1595 => x"74206661",
  1596 => x"696c6564",
  1597 => x"210a0000",
  1598 => x"53444843",
  1599 => x"20657272",
  1600 => x"6f72210a",
  1601 => x"00000000",
  1602 => x"57726974",
  1603 => x"65206661",
  1604 => x"696c6564",
  1605 => x"0a000000",
  1606 => x"52656164",
  1607 => x"20666169",
  1608 => x"6c65640a",
  1609 => x"00000000",
  1610 => x"43617264",
  1611 => x"20696e69",
  1612 => x"74206661",
  1613 => x"696c6564",
  1614 => x"0a000000",
  1615 => x"46415431",
  1616 => x"36202020",
  1617 => x"00000000",
  1618 => x"46415433",
  1619 => x"32202020",
  1620 => x"00000000",
  1621 => x"4e6f2070",
  1622 => x"61727469",
  1623 => x"74696f6e",
  1624 => x"20736967",
  1625 => x"0a000000",
  1626 => x"42616420",
  1627 => x"70617274",
  1628 => x"0a000000",
  1629 => x"4261636b",
  1630 => x"00000000",
  1631 => x"00000002",
  1632 => x"00000002",
  1633 => x"000017b0",
  1634 => x"00000000",
  1635 => x"00000002",
  1636 => x"000017c8",
  1637 => x"00000000",
  1638 => x"00000002",
  1639 => x"000017e0",
  1640 => x"0000034e",
  1641 => x"00000003",
  1642 => x"00001a24",
  1643 => x"00000004",
  1644 => x"00000003",
  1645 => x"00001a1c",
  1646 => x"00000002",
  1647 => x"00000003",
  1648 => x"00001a14",
  1649 => x"00000002",
  1650 => x"00000003",
  1651 => x"00001a0c",
  1652 => x"00000002",
  1653 => x"00000003",
  1654 => x"00001a04",
  1655 => x"00000002",
  1656 => x"00000002",
  1657 => x"000017e8",
  1658 => x"0000177b",
  1659 => x"00000002",
  1660 => x"00001800",
  1661 => x"000006bf",
  1662 => x"00000000",
  1663 => x"00000000",
  1664 => x"00000000",
  1665 => x"00001808",
  1666 => x"00001814",
  1667 => x"00001820",
  1668 => x"00001828",
  1669 => x"0000182c",
  1670 => x"0000183c",
  1671 => x"0000184c",
  1672 => x"0000185c",
  1673 => x"00001868",
  1674 => x"00001878",
  1675 => x"0000188c",
  1676 => x"000018a0",
  1677 => x"00000004",
  1678 => x"000018b4",
  1679 => x"00001a34",
  1680 => x"00000004",
  1681 => x"000018c4",
  1682 => x"00001980",
  1683 => x"00000000",
  1684 => x"00000000",
  1685 => x"00000000",
  1686 => x"00000000",
  1687 => x"00000000",
  1688 => x"00000000",
  1689 => x"00000000",
  1690 => x"00000000",
  1691 => x"00000000",
  1692 => x"00000000",
  1693 => x"00000000",
  1694 => x"00000000",
  1695 => x"00000000",
  1696 => x"00000000",
  1697 => x"00000000",
  1698 => x"00000000",
  1699 => x"00000000",
  1700 => x"00000000",
  1701 => x"00000000",
  1702 => x"00000000",
  1703 => x"00000000",
  1704 => x"00000000",
  1705 => x"00000000",
  1706 => x"00000000",
  1707 => x"00000002",
  1708 => x"00001f0c",
  1709 => x"0000157d",
  1710 => x"00000002",
  1711 => x"00001f2a",
  1712 => x"0000157d",
  1713 => x"00000002",
  1714 => x"00001f48",
  1715 => x"0000157d",
  1716 => x"00000002",
  1717 => x"00001f66",
  1718 => x"0000157d",
  1719 => x"00000002",
  1720 => x"00001f84",
  1721 => x"0000157d",
  1722 => x"00000002",
  1723 => x"00001fa2",
  1724 => x"0000157d",
  1725 => x"00000002",
  1726 => x"00001fc0",
  1727 => x"0000157d",
  1728 => x"00000002",
  1729 => x"00001fde",
  1730 => x"0000157d",
  1731 => x"00000002",
  1732 => x"00001ffc",
  1733 => x"0000157d",
  1734 => x"00000002",
  1735 => x"0000201a",
  1736 => x"0000157d",
  1737 => x"00000002",
  1738 => x"00002038",
  1739 => x"0000157d",
  1740 => x"00000002",
  1741 => x"00002056",
  1742 => x"0000157d",
  1743 => x"00000002",
  1744 => x"00002074",
  1745 => x"0000157d",
  1746 => x"00000004",
  1747 => x"00001974",
  1748 => x"00000000",
  1749 => x"00000000",
  1750 => x"00000000",
  1751 => x"0000170f",
  1752 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

